
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    ram_cell[       0] = 32'h00000037;
    ram_cell[       1] = 32'h000000a6;
    ram_cell[       2] = 32'h00000106;
    ram_cell[       3] = 32'h00000070;
    ram_cell[       4] = 32'h00000182;
    ram_cell[       5] = 32'h00000178;
    ram_cell[       6] = 32'h00000191;
    ram_cell[       7] = 32'h0000009f;
    ram_cell[       8] = 32'h000001e6;
    ram_cell[       9] = 32'h000000f6;
    ram_cell[      10] = 32'h0000012f;
    ram_cell[      11] = 32'h00000143;
    ram_cell[      12] = 32'h000000b0;
    ram_cell[      13] = 32'h00000114;
    ram_cell[      14] = 32'h00000102;
    ram_cell[      15] = 32'h000000ba;
    ram_cell[      16] = 32'h000001a6;
    ram_cell[      17] = 32'h000000b3;
    ram_cell[      18] = 32'h00000006;
    ram_cell[      19] = 32'h00000079;
    ram_cell[      20] = 32'h00000032;
    ram_cell[      21] = 32'h000001d0;
    ram_cell[      22] = 32'h000000e6;
    ram_cell[      23] = 32'h00000001;
    ram_cell[      24] = 32'h000001e2;
    ram_cell[      25] = 32'h000001f3;
    ram_cell[      26] = 32'h00000128;
    ram_cell[      27] = 32'h0000009e;
    ram_cell[      28] = 32'h0000010b;
    ram_cell[      29] = 32'h000001bf;
    ram_cell[      30] = 32'h000000b8;
    ram_cell[      31] = 32'h00000140;
    ram_cell[      32] = 32'h000000fd;
    ram_cell[      33] = 32'h000001f9;
    ram_cell[      34] = 32'h000001ad;
    ram_cell[      35] = 32'h00000003;
    ram_cell[      36] = 32'h000000e5;
    ram_cell[      37] = 32'h000001f2;
    ram_cell[      38] = 32'h000001d9;
    ram_cell[      39] = 32'h000000fb;
    ram_cell[      40] = 32'h00000199;
    ram_cell[      41] = 32'h000001e8;
    ram_cell[      42] = 32'h00000029;
    ram_cell[      43] = 32'h00000179;
    ram_cell[      44] = 32'h00000048;
    ram_cell[      45] = 32'h000000ab;
    ram_cell[      46] = 32'h000000ca;
    ram_cell[      47] = 32'h00000092;
    ram_cell[      48] = 32'h000001b3;
    ram_cell[      49] = 32'h000000a8;
    ram_cell[      50] = 32'h000001b9;
    ram_cell[      51] = 32'h000001f6;
    ram_cell[      52] = 32'h000001db;
    ram_cell[      53] = 32'h00000087;
    ram_cell[      54] = 32'h00000163;
    ram_cell[      55] = 32'h000001b0;
    ram_cell[      56] = 32'h00000185;
    ram_cell[      57] = 32'h000001af;
    ram_cell[      58] = 32'h000001c9;
    ram_cell[      59] = 32'h00000148;
    ram_cell[      60] = 32'h0000018f;
    ram_cell[      61] = 32'h00000186;
    ram_cell[      62] = 32'h0000001f;
    ram_cell[      63] = 32'h0000003c;
    ram_cell[      64] = 32'h00000142;
    ram_cell[      65] = 32'h00000164;
    ram_cell[      66] = 32'h0000014e;
    ram_cell[      67] = 32'h000000af;
    ram_cell[      68] = 32'h00000097;
    ram_cell[      69] = 32'h000001c0;
    ram_cell[      70] = 32'h0000017f;
    ram_cell[      71] = 32'h00000175;
    ram_cell[      72] = 32'h00000165;
    ram_cell[      73] = 32'h00000138;
    ram_cell[      74] = 32'h000001de;
    ram_cell[      75] = 32'h0000000c;
    ram_cell[      76] = 32'h00000065;
    ram_cell[      77] = 32'h00000085;
    ram_cell[      78] = 32'h00000031;
    ram_cell[      79] = 32'h0000016d;
    ram_cell[      80] = 32'h00000012;
    ram_cell[      81] = 32'h0000004a;
    ram_cell[      82] = 32'h00000055;
    ram_cell[      83] = 32'h000000f7;
    ram_cell[      84] = 32'h00000141;
    ram_cell[      85] = 32'h00000107;
    ram_cell[      86] = 32'h00000112;
    ram_cell[      87] = 32'h000001f5;
    ram_cell[      88] = 32'h000001d1;
    ram_cell[      89] = 32'h0000006f;
    ram_cell[      90] = 32'h0000016a;
    ram_cell[      91] = 32'h000000db;
    ram_cell[      92] = 32'h0000015c;
    ram_cell[      93] = 32'h0000000b;
    ram_cell[      94] = 32'h000001ca;
    ram_cell[      95] = 32'h00000062;
    ram_cell[      96] = 32'h00000159;
    ram_cell[      97] = 32'h00000197;
    ram_cell[      98] = 32'h0000015f;
    ram_cell[      99] = 32'h000001b4;
    ram_cell[     100] = 32'h00000093;
    ram_cell[     101] = 32'h000001e9;
    ram_cell[     102] = 32'h000000a9;
    ram_cell[     103] = 32'h00000111;
    ram_cell[     104] = 32'h000001a8;
    ram_cell[     105] = 32'h000000fa;
    ram_cell[     106] = 32'h0000004e;
    ram_cell[     107] = 32'h000000b6;
    ram_cell[     108] = 32'h000000c2;
    ram_cell[     109] = 32'h000001ed;
    ram_cell[     110] = 32'h0000000e;
    ram_cell[     111] = 32'h00000103;
    ram_cell[     112] = 32'h00000082;
    ram_cell[     113] = 32'h00000162;
    ram_cell[     114] = 32'h000000ce;
    ram_cell[     115] = 32'h00000124;
    ram_cell[     116] = 32'h00000115;
    ram_cell[     117] = 32'h000000df;
    ram_cell[     118] = 32'h000000e3;
    ram_cell[     119] = 32'h0000012e;
    ram_cell[     120] = 32'h000001c3;
    ram_cell[     121] = 32'h000001c7;
    ram_cell[     122] = 32'h000001ac;
    ram_cell[     123] = 32'h00000026;
    ram_cell[     124] = 32'h0000004c;
    ram_cell[     125] = 32'h00000108;
    ram_cell[     126] = 32'h00000060;
    ram_cell[     127] = 32'h000000bb;
    ram_cell[     128] = 32'h0000009c;
    ram_cell[     129] = 32'h00000068;
    ram_cell[     130] = 32'h00000033;
    ram_cell[     131] = 32'h0000015e;
    ram_cell[     132] = 32'h000000f5;
    ram_cell[     133] = 32'h00000195;
    ram_cell[     134] = 32'h00000025;
    ram_cell[     135] = 32'h00000018;
    ram_cell[     136] = 32'h0000006b;
    ram_cell[     137] = 32'h000001a5;
    ram_cell[     138] = 32'h00000147;
    ram_cell[     139] = 32'h00000189;
    ram_cell[     140] = 32'h00000132;
    ram_cell[     141] = 32'h00000027;
    ram_cell[     142] = 32'h00000135;
    ram_cell[     143] = 32'h0000019d;
    ram_cell[     144] = 32'h0000010a;
    ram_cell[     145] = 32'h000000ee;
    ram_cell[     146] = 32'h0000016b;
    ram_cell[     147] = 32'h00000158;
    ram_cell[     148] = 32'h000001f8;
    ram_cell[     149] = 32'h00000109;
    ram_cell[     150] = 32'h00000042;
    ram_cell[     151] = 32'h0000002e;
    ram_cell[     152] = 32'h00000083;
    ram_cell[     153] = 32'h00000020;
    ram_cell[     154] = 32'h000001bb;
    ram_cell[     155] = 32'h000000a4;
    ram_cell[     156] = 32'h000001e3;
    ram_cell[     157] = 32'h0000001c;
    ram_cell[     158] = 32'h0000004b;
    ram_cell[     159] = 32'h00000166;
    ram_cell[     160] = 32'h00000056;
    ram_cell[     161] = 32'h00000136;
    ram_cell[     162] = 32'h0000005c;
    ram_cell[     163] = 32'h00000067;
    ram_cell[     164] = 32'h00000170;
    ram_cell[     165] = 32'h000000eb;
    ram_cell[     166] = 32'h000000d1;
    ram_cell[     167] = 32'h00000014;
    ram_cell[     168] = 32'h0000019e;
    ram_cell[     169] = 32'h0000012a;
    ram_cell[     170] = 32'h000001ae;
    ram_cell[     171] = 32'h00000156;
    ram_cell[     172] = 32'h0000018c;
    ram_cell[     173] = 32'h00000155;
    ram_cell[     174] = 32'h0000011a;
    ram_cell[     175] = 32'h0000014d;
    ram_cell[     176] = 32'h000000b9;
    ram_cell[     177] = 32'h00000193;
    ram_cell[     178] = 32'h0000000d;
    ram_cell[     179] = 32'h000001cd;
    ram_cell[     180] = 32'h00000154;
    ram_cell[     181] = 32'h000000d5;
    ram_cell[     182] = 32'h000001b2;
    ram_cell[     183] = 32'h00000044;
    ram_cell[     184] = 32'h00000078;
    ram_cell[     185] = 32'h00000061;
    ram_cell[     186] = 32'h00000050;
    ram_cell[     187] = 32'h00000054;
    ram_cell[     188] = 32'h000001e7;
    ram_cell[     189] = 32'h0000005e;
    ram_cell[     190] = 32'h0000018a;
    ram_cell[     191] = 32'h00000121;
    ram_cell[     192] = 32'h00000075;
    ram_cell[     193] = 32'h000000c5;
    ram_cell[     194] = 32'h0000008d;
    ram_cell[     195] = 32'h000000ea;
    ram_cell[     196] = 32'h00000180;
    ram_cell[     197] = 32'h000000b7;
    ram_cell[     198] = 32'h000000d7;
    ram_cell[     199] = 32'h0000002c;
    ram_cell[     200] = 32'h000000ae;
    ram_cell[     201] = 32'h000001c1;
    ram_cell[     202] = 32'h000000ed;
    ram_cell[     203] = 32'h0000018e;
    ram_cell[     204] = 32'h00000118;
    ram_cell[     205] = 32'h000001e5;
    ram_cell[     206] = 32'h000001ea;
    ram_cell[     207] = 32'h00000011;
    ram_cell[     208] = 32'h000001d2;
    ram_cell[     209] = 32'h00000119;
    ram_cell[     210] = 32'h0000015d;
    ram_cell[     211] = 32'h00000113;
    ram_cell[     212] = 32'h00000059;
    ram_cell[     213] = 32'h000000cc;
    ram_cell[     214] = 32'h000000d4;
    ram_cell[     215] = 32'h00000110;
    ram_cell[     216] = 32'h00000015;
    ram_cell[     217] = 32'h000000ec;
    ram_cell[     218] = 32'h00000122;
    ram_cell[     219] = 32'h00000051;
    ram_cell[     220] = 32'h000001aa;
    ram_cell[     221] = 32'h00000120;
    ram_cell[     222] = 32'h00000072;
    ram_cell[     223] = 32'h000001ef;
    ram_cell[     224] = 32'h00000081;
    ram_cell[     225] = 32'h000000f9;
    ram_cell[     226] = 32'h0000014f;
    ram_cell[     227] = 32'h000001fc;
    ram_cell[     228] = 32'h000000c7;
    ram_cell[     229] = 32'h0000006c;
    ram_cell[     230] = 32'h0000007a;
    ram_cell[     231] = 32'h0000009b;
    ram_cell[     232] = 32'h0000019a;
    ram_cell[     233] = 32'h00000047;
    ram_cell[     234] = 32'h000001e0;
    ram_cell[     235] = 32'h00000137;
    ram_cell[     236] = 32'h00000004;
    ram_cell[     237] = 32'h0000002f;
    ram_cell[     238] = 32'h0000016f;
    ram_cell[     239] = 32'h000000bd;
    ram_cell[     240] = 32'h00000035;
    ram_cell[     241] = 32'h000001df;
    ram_cell[     242] = 32'h0000007e;
    ram_cell[     243] = 32'h00000000;
    ram_cell[     244] = 32'h00000038;
    ram_cell[     245] = 32'h00000016;
    ram_cell[     246] = 32'h0000011f;
    ram_cell[     247] = 32'h00000160;
    ram_cell[     248] = 32'h000001a1;
    ram_cell[     249] = 32'h00000100;
    ram_cell[     250] = 32'h000000b5;
    ram_cell[     251] = 32'h000001eb;
    ram_cell[     252] = 32'h00000058;
    ram_cell[     253] = 32'h000000e7;
    ram_cell[     254] = 32'h0000019f;
    ram_cell[     255] = 32'h00000049;
    ram_cell[     256] = 32'h0000001d;
    ram_cell[     257] = 32'h0000000f;
    ram_cell[     258] = 32'h000001f0;
    ram_cell[     259] = 32'h0000003e;
    ram_cell[     260] = 32'h000000e8;
    ram_cell[     261] = 32'h000000cf;
    ram_cell[     262] = 32'h00000144;
    ram_cell[     263] = 32'h00000019;
    ram_cell[     264] = 32'h00000125;
    ram_cell[     265] = 32'h000001a7;
    ram_cell[     266] = 32'h0000012d;
    ram_cell[     267] = 32'h0000013f;
    ram_cell[     268] = 32'h0000013d;
    ram_cell[     269] = 32'h000000ac;
    ram_cell[     270] = 32'h00000017;
    ram_cell[     271] = 32'h000001c8;
    ram_cell[     272] = 32'h00000030;
    ram_cell[     273] = 32'h0000004f;
    ram_cell[     274] = 32'h00000150;
    ram_cell[     275] = 32'h000000f8;
    ram_cell[     276] = 32'h000001c6;
    ram_cell[     277] = 32'h000000d8;
    ram_cell[     278] = 32'h0000002a;
    ram_cell[     279] = 32'h0000013e;
    ram_cell[     280] = 32'h0000008f;
    ram_cell[     281] = 32'h000000ff;
    ram_cell[     282] = 32'h000001fb;
    ram_cell[     283] = 32'h00000021;
    ram_cell[     284] = 32'h00000133;
    ram_cell[     285] = 32'h0000014b;
    ram_cell[     286] = 32'h000001a4;
    ram_cell[     287] = 32'h00000126;
    ram_cell[     288] = 32'h0000013b;
    ram_cell[     289] = 32'h0000015a;
    ram_cell[     290] = 32'h000001ba;
    ram_cell[     291] = 32'h0000012c;
    ram_cell[     292] = 32'h000001f1;
    ram_cell[     293] = 32'h000000bf;
    ram_cell[     294] = 32'h00000066;
    ram_cell[     295] = 32'h0000008b;
    ram_cell[     296] = 32'h000000f2;
    ram_cell[     297] = 32'h00000183;
    ram_cell[     298] = 32'h000001c5;
    ram_cell[     299] = 32'h00000077;
    ram_cell[     300] = 32'h000001ab;
    ram_cell[     301] = 32'h0000001e;
    ram_cell[     302] = 32'h000000a5;
    ram_cell[     303] = 32'h00000190;
    ram_cell[     304] = 32'h00000034;
    ram_cell[     305] = 32'h00000173;
    ram_cell[     306] = 32'h0000004d;
    ram_cell[     307] = 32'h0000008c;
    ram_cell[     308] = 32'h000001d8;
    ram_cell[     309] = 32'h00000052;
    ram_cell[     310] = 32'h000001c2;
    ram_cell[     311] = 32'h0000018b;
    ram_cell[     312] = 32'h00000098;
    ram_cell[     313] = 32'h000000b1;
    ram_cell[     314] = 32'h00000167;
    ram_cell[     315] = 32'h0000017b;
    ram_cell[     316] = 32'h000000d0;
    ram_cell[     317] = 32'h00000053;
    ram_cell[     318] = 32'h00000073;
    ram_cell[     319] = 32'h000000f3;
    ram_cell[     320] = 32'h0000011e;
    ram_cell[     321] = 32'h0000003a;
    ram_cell[     322] = 32'h00000194;
    ram_cell[     323] = 32'h00000131;
    ram_cell[     324] = 32'h00000010;
    ram_cell[     325] = 32'h000000b2;
    ram_cell[     326] = 32'h0000002b;
    ram_cell[     327] = 32'h0000010d;
    ram_cell[     328] = 32'h00000151;
    ram_cell[     329] = 32'h00000184;
    ram_cell[     330] = 32'h0000010e;
    ram_cell[     331] = 32'h000001c4;
    ram_cell[     332] = 32'h000001cc;
    ram_cell[     333] = 32'h0000013c;
    ram_cell[     334] = 32'h0000001b;
    ram_cell[     335] = 32'h00000104;
    ram_cell[     336] = 32'h00000074;
    ram_cell[     337] = 32'h00000089;
    ram_cell[     338] = 32'h0000015b;
    ram_cell[     339] = 32'h00000196;
    ram_cell[     340] = 32'h00000009;
    ram_cell[     341] = 32'h000000cd;
    ram_cell[     342] = 32'h00000134;
    ram_cell[     343] = 32'h000000aa;
    ram_cell[     344] = 32'h000000dc;
    ram_cell[     345] = 32'h000001cb;
    ram_cell[     346] = 32'h000001b7;
    ram_cell[     347] = 32'h0000005b;
    ram_cell[     348] = 32'h00000172;
    ram_cell[     349] = 32'h00000091;
    ram_cell[     350] = 32'h00000116;
    ram_cell[     351] = 32'h00000071;
    ram_cell[     352] = 32'h00000168;
    ram_cell[     353] = 32'h00000105;
    ram_cell[     354] = 32'h00000036;
    ram_cell[     355] = 32'h000001fa;
    ram_cell[     356] = 32'h00000174;
    ram_cell[     357] = 32'h000000dd;
    ram_cell[     358] = 32'h000001d7;
    ram_cell[     359] = 32'h000000d9;
    ram_cell[     360] = 32'h000000c9;
    ram_cell[     361] = 32'h000001ff;
    ram_cell[     362] = 32'h0000005d;
    ram_cell[     363] = 32'h0000018d;
    ram_cell[     364] = 32'h00000171;
    ram_cell[     365] = 32'h0000008a;
    ram_cell[     366] = 32'h0000017c;
    ram_cell[     367] = 32'h000000d2;
    ram_cell[     368] = 32'h000000c4;
    ram_cell[     369] = 32'h00000084;
    ram_cell[     370] = 32'h00000022;
    ram_cell[     371] = 32'h00000149;
    ram_cell[     372] = 32'h0000005a;
    ram_cell[     373] = 32'h00000094;
    ram_cell[     374] = 32'h000001bc;
    ram_cell[     375] = 32'h000000c3;
    ram_cell[     376] = 32'h00000145;
    ram_cell[     377] = 32'h000000c1;
    ram_cell[     378] = 32'h0000000a;
    ram_cell[     379] = 32'h000001fe;
    ram_cell[     380] = 32'h000000be;
    ram_cell[     381] = 32'h000001ec;
    ram_cell[     382] = 32'h000000f4;
    ram_cell[     383] = 32'h0000003d;
    ram_cell[     384] = 32'h00000039;
    ram_cell[     385] = 32'h00000088;
    ram_cell[     386] = 32'h00000076;
    ram_cell[     387] = 32'h00000045;
    ram_cell[     388] = 32'h000000c0;
    ram_cell[     389] = 32'h000000fc;
    ram_cell[     390] = 32'h000001a0;
    ram_cell[     391] = 32'h00000192;
    ram_cell[     392] = 32'h00000063;
    ram_cell[     393] = 32'h000001d5;
    ram_cell[     394] = 32'h00000005;
    ram_cell[     395] = 32'h000001a3;
    ram_cell[     396] = 32'h0000002d;
    ram_cell[     397] = 32'h0000019b;
    ram_cell[     398] = 32'h000001b8;
    ram_cell[     399] = 32'h000000c6;
    ram_cell[     400] = 32'h000000bc;
    ram_cell[     401] = 32'h000001bd;
    ram_cell[     402] = 32'h0000017e;
    ram_cell[     403] = 32'h0000014a;
    ram_cell[     404] = 32'h00000069;
    ram_cell[     405] = 32'h000001b1;
    ram_cell[     406] = 32'h00000101;
    ram_cell[     407] = 32'h0000010f;
    ram_cell[     408] = 32'h00000057;
    ram_cell[     409] = 32'h000001b5;
    ram_cell[     410] = 32'h00000127;
    ram_cell[     411] = 32'h00000187;
    ram_cell[     412] = 32'h00000086;
    ram_cell[     413] = 32'h0000006e;
    ram_cell[     414] = 32'h0000007d;
    ram_cell[     415] = 32'h00000198;
    ram_cell[     416] = 32'h000001b6;
    ram_cell[     417] = 32'h00000024;
    ram_cell[     418] = 32'h0000009a;
    ram_cell[     419] = 32'h000001a9;
    ram_cell[     420] = 32'h00000064;
    ram_cell[     421] = 32'h0000003f;
    ram_cell[     422] = 32'h0000011b;
    ram_cell[     423] = 32'h000001a2;
    ram_cell[     424] = 32'h0000019c;
    ram_cell[     425] = 32'h00000157;
    ram_cell[     426] = 32'h00000043;
    ram_cell[     427] = 32'h000000ef;
    ram_cell[     428] = 32'h00000040;
    ram_cell[     429] = 32'h0000003b;
    ram_cell[     430] = 32'h000000f0;
    ram_cell[     431] = 32'h000001d6;
    ram_cell[     432] = 32'h0000016c;
    ram_cell[     433] = 32'h00000028;
    ram_cell[     434] = 32'h000000a7;
    ram_cell[     435] = 32'h00000169;
    ram_cell[     436] = 32'h000001dd;
    ram_cell[     437] = 32'h0000007f;
    ram_cell[     438] = 32'h000000d3;
    ram_cell[     439] = 32'h0000012b;
    ram_cell[     440] = 32'h0000001a;
    ram_cell[     441] = 32'h000000cb;
    ram_cell[     442] = 32'h00000046;
    ram_cell[     443] = 32'h000000a2;
    ram_cell[     444] = 32'h000001dc;
    ram_cell[     445] = 32'h0000009d;
    ram_cell[     446] = 32'h000000fe;
    ram_cell[     447] = 32'h000000a1;
    ram_cell[     448] = 32'h000001d3;
    ram_cell[     449] = 32'h000000a3;
    ram_cell[     450] = 32'h00000161;
    ram_cell[     451] = 32'h000000de;
    ram_cell[     452] = 32'h00000188;
    ram_cell[     453] = 32'h000001f7;
    ram_cell[     454] = 32'h00000152;
    ram_cell[     455] = 32'h00000139;
    ram_cell[     456] = 32'h0000007c;
    ram_cell[     457] = 32'h00000023;
    ram_cell[     458] = 32'h0000013a;
    ram_cell[     459] = 32'h000001cf;
    ram_cell[     460] = 32'h000001ee;
    ram_cell[     461] = 32'h00000146;
    ram_cell[     462] = 32'h000000d6;
    ram_cell[     463] = 32'h00000153;
    ram_cell[     464] = 32'h000000da;
    ram_cell[     465] = 32'h000001d4;
    ram_cell[     466] = 32'h0000007b;
    ram_cell[     467] = 32'h00000080;
    ram_cell[     468] = 32'h000000e2;
    ram_cell[     469] = 32'h000000e4;
    ram_cell[     470] = 32'h00000007;
    ram_cell[     471] = 32'h00000095;
    ram_cell[     472] = 32'h0000016e;
    ram_cell[     473] = 32'h000000b4;
    ram_cell[     474] = 32'h00000090;
    ram_cell[     475] = 32'h0000014c;
    ram_cell[     476] = 32'h00000002;
    ram_cell[     477] = 32'h000000e0;
    ram_cell[     478] = 32'h000000c8;
    ram_cell[     479] = 32'h0000011c;
    ram_cell[     480] = 32'h00000008;
    ram_cell[     481] = 32'h0000006a;
    ram_cell[     482] = 32'h00000176;
    ram_cell[     483] = 32'h0000011d;
    ram_cell[     484] = 32'h000001e4;
    ram_cell[     485] = 32'h000001da;
    ram_cell[     486] = 32'h0000017a;
    ram_cell[     487] = 32'h000001e1;
    ram_cell[     488] = 32'h0000006d;
    ram_cell[     489] = 32'h00000013;
    ram_cell[     490] = 32'h000000e9;
    ram_cell[     491] = 32'h00000117;
    ram_cell[     492] = 32'h000001f4;
    ram_cell[     493] = 32'h00000177;
    ram_cell[     494] = 32'h0000005f;
    ram_cell[     495] = 32'h00000130;
    ram_cell[     496] = 32'h000000a0;
    ram_cell[     497] = 32'h000000e1;
    ram_cell[     498] = 32'h00000129;
    ram_cell[     499] = 32'h000000f1;
    ram_cell[     500] = 32'h0000017d;
    ram_cell[     501] = 32'h0000010c;
    ram_cell[     502] = 32'h000001fd;
    ram_cell[     503] = 32'h000000ad;
    ram_cell[     504] = 32'h0000008e;
    ram_cell[     505] = 32'h000001ce;
    ram_cell[     506] = 32'h00000123;
    ram_cell[     507] = 32'h00000099;
    ram_cell[     508] = 32'h000001be;
    ram_cell[     509] = 32'h00000096;
    ram_cell[     510] = 32'h00000041;
    ram_cell[     511] = 32'h00000181;
end

endmodule




// module mem #(                   // 
// parameter  ADDR_LEN  = 11   // 
// ) (
// input  clk, rst,
// input  [ADDR_LEN-1:0] addr, // memory address
// output reg [31:0] rd_data,  // data read out
// input  wr_req,
// input  [31:0] wr_data       // data write in
// );
// localparam MEM_SIZE = 1<<ADDR_LEN;
// reg [31:0] ram_cell [MEM_SIZE];

// always @ (posedge clk or posedge rst)
// if(rst)
//     rd_data <= 0;
// else
//     rd_data <= ram_cell[addr];

// always @ (posedge clk)
// if(wr_req) 
//     ram_cell[addr] <= wr_data;

// initial begin
// // dst matrix C
// ram_cell[       0] = 32'h0;  // 32'h3c58db17;
// ram_cell[       1] = 32'h0;  // 32'h94e418a6;
// ram_cell[       2] = 32'h0;  // 32'h09f9452d;
// ram_cell[       3] = 32'h0;  // 32'h81b8aa66;
// ram_cell[       4] = 32'h0;  // 32'h9adcdee3;
// ram_cell[       5] = 32'h0;  // 32'hf809994c;
// ram_cell[       6] = 32'h0;  // 32'ha1ca7f52;
// ram_cell[       7] = 32'h0;  // 32'h2f76e1d1;
// ram_cell[       8] = 32'h0;  // 32'h641e4889;
// ram_cell[       9] = 32'h0;  // 32'hd24b35cd;
// ram_cell[      10] = 32'h0;  // 32'hc9db24f7;
// ram_cell[      11] = 32'h0;  // 32'hc33f8da3;
// ram_cell[      12] = 32'h0;  // 32'hd6cdad70;
// ram_cell[      13] = 32'h0;  // 32'h2f9906ff;
// ram_cell[      14] = 32'h0;  // 32'haaa78bc8;
// ram_cell[      15] = 32'h0;  // 32'h678bcbcd;
// ram_cell[      16] = 32'h0;  // 32'h6f925258;
// ram_cell[      17] = 32'h0;  // 32'h1350f68c;
// ram_cell[      18] = 32'h0;  // 32'h61004b31;
// ram_cell[      19] = 32'h0;  // 32'h9672dc82;
// ram_cell[      20] = 32'h0;  // 32'h724b8521;
// ram_cell[      21] = 32'h0;  // 32'ha27c51c8;
// ram_cell[      22] = 32'h0;  // 32'h9dc4128a;
// ram_cell[      23] = 32'h0;  // 32'h24d0160a;
// ram_cell[      24] = 32'h0;  // 32'h5b3f0dd9;
// ram_cell[      25] = 32'h0;  // 32'hef9ffd28;
// ram_cell[      26] = 32'h0;  // 32'hfa600d55;
// ram_cell[      27] = 32'h0;  // 32'h8c593f82;
// ram_cell[      28] = 32'h0;  // 32'h1994d141;
// ram_cell[      29] = 32'h0;  // 32'h8c92456c;
// ram_cell[      30] = 32'h0;  // 32'h7be5d474;
// ram_cell[      31] = 32'h0;  // 32'hd9181b06;
// ram_cell[      32] = 32'h0;  // 32'hbf2a0b2e;
// ram_cell[      33] = 32'h0;  // 32'hc0438cc5;
// ram_cell[      34] = 32'h0;  // 32'hd9ee0b1b;
// ram_cell[      35] = 32'h0;  // 32'h4d805b2c;
// ram_cell[      36] = 32'h0;  // 32'h5ff1f603;
// ram_cell[      37] = 32'h0;  // 32'h9bcd04d2;
// ram_cell[      38] = 32'h0;  // 32'h4ad235ab;
// ram_cell[      39] = 32'h0;  // 32'h00edeef2;
// ram_cell[      40] = 32'h0;  // 32'h2d04801c;
// ram_cell[      41] = 32'h0;  // 32'h42551ff3;
// ram_cell[      42] = 32'h0;  // 32'hbb5ed37b;
// ram_cell[      43] = 32'h0;  // 32'hfd0e61f3;
// ram_cell[      44] = 32'h0;  // 32'h42fe10b5;
// ram_cell[      45] = 32'h0;  // 32'h56b31c0f;
// ram_cell[      46] = 32'h0;  // 32'h6a0a2983;
// ram_cell[      47] = 32'h0;  // 32'h839d0d5b;
// ram_cell[      48] = 32'h0;  // 32'h3a7933a2;
// ram_cell[      49] = 32'h0;  // 32'h943e7942;
// ram_cell[      50] = 32'h0;  // 32'h71dcfc65;
// ram_cell[      51] = 32'h0;  // 32'h2a812803;
// ram_cell[      52] = 32'h0;  // 32'h7b33e05a;
// ram_cell[      53] = 32'h0;  // 32'h7ddb6cbb;
// ram_cell[      54] = 32'h0;  // 32'h77eb6a7a;
// ram_cell[      55] = 32'h0;  // 32'h2ffabf86;
// ram_cell[      56] = 32'h0;  // 32'hbae41542;
// ram_cell[      57] = 32'h0;  // 32'h36013d95;
// ram_cell[      58] = 32'h0;  // 32'hf21d8c79;
// ram_cell[      59] = 32'h0;  // 32'he2c2f383;
// ram_cell[      60] = 32'h0;  // 32'h893f9c39;
// ram_cell[      61] = 32'h0;  // 32'h50d86d3b;
// ram_cell[      62] = 32'h0;  // 32'h17aa3945;
// ram_cell[      63] = 32'h0;  // 32'h42dc5eb4;
// ram_cell[      64] = 32'h0;  // 32'h69f9d176;
// ram_cell[      65] = 32'h0;  // 32'hb5caf8a0;
// ram_cell[      66] = 32'h0;  // 32'h0f32c73e;
// ram_cell[      67] = 32'h0;  // 32'hc5dc6696;
// ram_cell[      68] = 32'h0;  // 32'h8267e53b;
// ram_cell[      69] = 32'h0;  // 32'h0bb15a0b;
// ram_cell[      70] = 32'h0;  // 32'h7b50a2f1;
// ram_cell[      71] = 32'h0;  // 32'h1f0380f9;
// ram_cell[      72] = 32'h0;  // 32'hccf587f7;
// ram_cell[      73] = 32'h0;  // 32'hb1b3bfa4;
// ram_cell[      74] = 32'h0;  // 32'h81939c5d;
// ram_cell[      75] = 32'h0;  // 32'h170b8766;
// ram_cell[      76] = 32'h0;  // 32'h9fc9345b;
// ram_cell[      77] = 32'h0;  // 32'h652d9631;
// ram_cell[      78] = 32'h0;  // 32'h7b75feba;
// ram_cell[      79] = 32'h0;  // 32'h8d5be980;
// ram_cell[      80] = 32'h0;  // 32'h121f4482;
// ram_cell[      81] = 32'h0;  // 32'h75bc24ce;
// ram_cell[      82] = 32'h0;  // 32'h391c5a3a;
// ram_cell[      83] = 32'h0;  // 32'h72dd99ac;
// ram_cell[      84] = 32'h0;  // 32'h9a3ac738;
// ram_cell[      85] = 32'h0;  // 32'h2bf863ef;
// ram_cell[      86] = 32'h0;  // 32'ha18c28b6;
// ram_cell[      87] = 32'h0;  // 32'h94559e38;
// ram_cell[      88] = 32'h0;  // 32'hd655b39b;
// ram_cell[      89] = 32'h0;  // 32'hedce726c;
// ram_cell[      90] = 32'h0;  // 32'h84b5da2b;
// ram_cell[      91] = 32'h0;  // 32'he4de3a06;
// ram_cell[      92] = 32'h0;  // 32'hc632a3be;
// ram_cell[      93] = 32'h0;  // 32'hcecd39d8;
// ram_cell[      94] = 32'h0;  // 32'ha882ac5b;
// ram_cell[      95] = 32'h0;  // 32'hdd1be2f4;
// ram_cell[      96] = 32'h0;  // 32'hb08b766b;
// ram_cell[      97] = 32'h0;  // 32'hc14931d9;
// ram_cell[      98] = 32'h0;  // 32'hdd1ff796;
// ram_cell[      99] = 32'h0;  // 32'h571c755f;
// ram_cell[     100] = 32'h0;  // 32'he4350195;
// ram_cell[     101] = 32'h0;  // 32'h3893aa35;
// ram_cell[     102] = 32'h0;  // 32'h15d6f84e;
// ram_cell[     103] = 32'h0;  // 32'h70f4dbf5;
// ram_cell[     104] = 32'h0;  // 32'hcf3152e5;
// ram_cell[     105] = 32'h0;  // 32'hbe910ff5;
// ram_cell[     106] = 32'h0;  // 32'h0d8ce6dd;
// ram_cell[     107] = 32'h0;  // 32'h71dec6bd;
// ram_cell[     108] = 32'h0;  // 32'hcb03d6d9;
// ram_cell[     109] = 32'h0;  // 32'h24282d91;
// ram_cell[     110] = 32'h0;  // 32'hb0bcdaaa;
// ram_cell[     111] = 32'h0;  // 32'h39eed65b;
// ram_cell[     112] = 32'h0;  // 32'h495da131;
// ram_cell[     113] = 32'h0;  // 32'hb271d4cd;
// ram_cell[     114] = 32'h0;  // 32'h7f2b37f3;
// ram_cell[     115] = 32'h0;  // 32'hf823bee0;
// ram_cell[     116] = 32'h0;  // 32'h0bcb7b98;
// ram_cell[     117] = 32'h0;  // 32'hbaf8cabd;
// ram_cell[     118] = 32'h0;  // 32'hda49c899;
// ram_cell[     119] = 32'h0;  // 32'h435a279b;
// ram_cell[     120] = 32'h0;  // 32'h6b775e98;
// ram_cell[     121] = 32'h0;  // 32'hf6fbfbaa;
// ram_cell[     122] = 32'h0;  // 32'hd9574182;
// ram_cell[     123] = 32'h0;  // 32'hd85452b4;
// ram_cell[     124] = 32'h0;  // 32'he897dd39;
// ram_cell[     125] = 32'h0;  // 32'h002588e5;
// ram_cell[     126] = 32'h0;  // 32'hfc0f7674;
// ram_cell[     127] = 32'h0;  // 32'h8a3ccbc2;
// ram_cell[     128] = 32'h0;  // 32'h783346a5;
// ram_cell[     129] = 32'h0;  // 32'h281ef16f;
// ram_cell[     130] = 32'h0;  // 32'h1b0bbf7a;
// ram_cell[     131] = 32'h0;  // 32'h44682b4c;
// ram_cell[     132] = 32'h0;  // 32'h7915b814;
// ram_cell[     133] = 32'h0;  // 32'he4c48b42;
// ram_cell[     134] = 32'h0;  // 32'h0df63eb3;
// ram_cell[     135] = 32'h0;  // 32'h7d919681;
// ram_cell[     136] = 32'h0;  // 32'hc6774295;
// ram_cell[     137] = 32'h0;  // 32'he85b4daa;
// ram_cell[     138] = 32'h0;  // 32'h55a3c5be;
// ram_cell[     139] = 32'h0;  // 32'h5b3f735c;
// ram_cell[     140] = 32'h0;  // 32'h3c1476c5;
// ram_cell[     141] = 32'h0;  // 32'h1cc9341e;
// ram_cell[     142] = 32'h0;  // 32'h56aebc60;
// ram_cell[     143] = 32'h0;  // 32'hde644135;
// ram_cell[     144] = 32'h0;  // 32'hc6dd3256;
// ram_cell[     145] = 32'h0;  // 32'hafd6be00;
// ram_cell[     146] = 32'h0;  // 32'hcda3ca02;
// ram_cell[     147] = 32'h0;  // 32'hda1b64b2;
// ram_cell[     148] = 32'h0;  // 32'h2cf59a79;
// ram_cell[     149] = 32'h0;  // 32'h6029fcf7;
// ram_cell[     150] = 32'h0;  // 32'he949abfd;
// ram_cell[     151] = 32'h0;  // 32'hc89498ad;
// ram_cell[     152] = 32'h0;  // 32'hace178c8;
// ram_cell[     153] = 32'h0;  // 32'hc9899839;
// ram_cell[     154] = 32'h0;  // 32'ha1527533;
// ram_cell[     155] = 32'h0;  // 32'he71dfba0;
// ram_cell[     156] = 32'h0;  // 32'hb4d42203;
// ram_cell[     157] = 32'h0;  // 32'h7259dd7c;
// ram_cell[     158] = 32'h0;  // 32'h96e04ce5;
// ram_cell[     159] = 32'h0;  // 32'h359cc056;
// ram_cell[     160] = 32'h0;  // 32'hb7a38799;
// ram_cell[     161] = 32'h0;  // 32'hed485009;
// ram_cell[     162] = 32'h0;  // 32'h2f5c0535;
// ram_cell[     163] = 32'h0;  // 32'h39d78498;
// ram_cell[     164] = 32'h0;  // 32'h770dcb44;
// ram_cell[     165] = 32'h0;  // 32'h5b300960;
// ram_cell[     166] = 32'h0;  // 32'h98d41d10;
// ram_cell[     167] = 32'h0;  // 32'h194e6ee6;
// ram_cell[     168] = 32'h0;  // 32'h6ca6a1e7;
// ram_cell[     169] = 32'h0;  // 32'hddd701c6;
// ram_cell[     170] = 32'h0;  // 32'h9086cd82;
// ram_cell[     171] = 32'h0;  // 32'h3698829e;
// ram_cell[     172] = 32'h0;  // 32'hfe3add20;
// ram_cell[     173] = 32'h0;  // 32'h213e964d;
// ram_cell[     174] = 32'h0;  // 32'ha1a4a1a4;
// ram_cell[     175] = 32'h0;  // 32'h2719dd9c;
// ram_cell[     176] = 32'h0;  // 32'hfd764f52;
// ram_cell[     177] = 32'h0;  // 32'h0c008ce8;
// ram_cell[     178] = 32'h0;  // 32'hf48b394c;
// ram_cell[     179] = 32'h0;  // 32'h622b5503;
// ram_cell[     180] = 32'h0;  // 32'h66896642;
// ram_cell[     181] = 32'h0;  // 32'ha3769d03;
// ram_cell[     182] = 32'h0;  // 32'h68057da1;
// ram_cell[     183] = 32'h0;  // 32'hfd8a3f6e;
// ram_cell[     184] = 32'h0;  // 32'h93b73e80;
// ram_cell[     185] = 32'h0;  // 32'hee182118;
// ram_cell[     186] = 32'h0;  // 32'h4c4b579e;
// ram_cell[     187] = 32'h0;  // 32'h292b8280;
// ram_cell[     188] = 32'h0;  // 32'h8bbaadd8;
// ram_cell[     189] = 32'h0;  // 32'hf0657406;
// ram_cell[     190] = 32'h0;  // 32'h2f2f7882;
// ram_cell[     191] = 32'h0;  // 32'hd7928396;
// ram_cell[     192] = 32'h0;  // 32'ha59e3068;
// ram_cell[     193] = 32'h0;  // 32'h743963cf;
// ram_cell[     194] = 32'h0;  // 32'habfcd4e8;
// ram_cell[     195] = 32'h0;  // 32'h206e68c0;
// ram_cell[     196] = 32'h0;  // 32'h8542c261;
// ram_cell[     197] = 32'h0;  // 32'h88e876c7;
// ram_cell[     198] = 32'h0;  // 32'h439645ff;
// ram_cell[     199] = 32'h0;  // 32'h6dd8912d;
// ram_cell[     200] = 32'h0;  // 32'h454729e9;
// ram_cell[     201] = 32'h0;  // 32'h046c3a50;
// ram_cell[     202] = 32'h0;  // 32'hfce4ee77;
// ram_cell[     203] = 32'h0;  // 32'h7170acbe;
// ram_cell[     204] = 32'h0;  // 32'hc870de7b;
// ram_cell[     205] = 32'h0;  // 32'h8e7af611;
// ram_cell[     206] = 32'h0;  // 32'h9f982dcb;
// ram_cell[     207] = 32'h0;  // 32'h006e6787;
// ram_cell[     208] = 32'h0;  // 32'hfc46fd59;
// ram_cell[     209] = 32'h0;  // 32'h43c982bb;
// ram_cell[     210] = 32'h0;  // 32'h52cfae64;
// ram_cell[     211] = 32'h0;  // 32'h85004632;
// ram_cell[     212] = 32'h0;  // 32'hc4d7672a;
// ram_cell[     213] = 32'h0;  // 32'h1130ed0c;
// ram_cell[     214] = 32'h0;  // 32'h3b15c773;
// ram_cell[     215] = 32'h0;  // 32'h229810d1;
// ram_cell[     216] = 32'h0;  // 32'h2f19594e;
// ram_cell[     217] = 32'h0;  // 32'h255359bd;
// ram_cell[     218] = 32'h0;  // 32'h45762ab2;
// ram_cell[     219] = 32'h0;  // 32'h09a08cd2;
// ram_cell[     220] = 32'h0;  // 32'h2ccfc44d;
// ram_cell[     221] = 32'h0;  // 32'h0033ad3b;
// ram_cell[     222] = 32'h0;  // 32'h4050afe4;
// ram_cell[     223] = 32'h0;  // 32'h5ad985e1;
// ram_cell[     224] = 32'h0;  // 32'hdcd042e1;
// ram_cell[     225] = 32'h0;  // 32'h39a49fd1;
// ram_cell[     226] = 32'h0;  // 32'h9564de5e;
// ram_cell[     227] = 32'h0;  // 32'h9c75fe89;
// ram_cell[     228] = 32'h0;  // 32'h51104768;
// ram_cell[     229] = 32'h0;  // 32'h44ba2a68;
// ram_cell[     230] = 32'h0;  // 32'hf022c7f4;
// ram_cell[     231] = 32'h0;  // 32'hfe7e594e;
// ram_cell[     232] = 32'h0;  // 32'h0c555151;
// ram_cell[     233] = 32'h0;  // 32'h4ba0a68f;
// ram_cell[     234] = 32'h0;  // 32'hb7021bab;
// ram_cell[     235] = 32'h0;  // 32'h99b49c5c;
// ram_cell[     236] = 32'h0;  // 32'h131c243e;
// ram_cell[     237] = 32'h0;  // 32'ha0df87d1;
// ram_cell[     238] = 32'h0;  // 32'h8247a3cf;
// ram_cell[     239] = 32'h0;  // 32'h6de3f215;
// ram_cell[     240] = 32'h0;  // 32'h646df1b5;
// ram_cell[     241] = 32'h0;  // 32'h560b4633;
// ram_cell[     242] = 32'h0;  // 32'h9bd255f6;
// ram_cell[     243] = 32'h0;  // 32'h446f4eb4;
// ram_cell[     244] = 32'h0;  // 32'h16c0bf76;
// ram_cell[     245] = 32'h0;  // 32'hd507cd24;
// ram_cell[     246] = 32'h0;  // 32'hbf14689e;
// ram_cell[     247] = 32'h0;  // 32'ha3ebd0f5;
// ram_cell[     248] = 32'h0;  // 32'h2897aea9;
// ram_cell[     249] = 32'h0;  // 32'h79c6eca7;
// ram_cell[     250] = 32'h0;  // 32'h88fb0f29;
// ram_cell[     251] = 32'h0;  // 32'h0875ee8a;
// ram_cell[     252] = 32'h0;  // 32'h0f85375d;
// ram_cell[     253] = 32'h0;  // 32'h2bcb9bac;
// ram_cell[     254] = 32'h0;  // 32'hc5ff889c;
// ram_cell[     255] = 32'h0;  // 32'hf4e8a784;
// // src matrix A
// ram_cell[     256] = 32'h67c69e3e;
// ram_cell[     257] = 32'ha45ad965;
// ram_cell[     258] = 32'hf9a5af28;
// ram_cell[     259] = 32'h96e488c5;
// ram_cell[     260] = 32'h8b369be4;
// ram_cell[     261] = 32'haaa89ec0;
// ram_cell[     262] = 32'h654875a4;
// ram_cell[     263] = 32'hd330fd7e;
// ram_cell[     264] = 32'h3b11ce13;
// ram_cell[     265] = 32'h760d6d22;
// ram_cell[     266] = 32'h80c41bf3;
// ram_cell[     267] = 32'hf00fdf20;
// ram_cell[     268] = 32'h208b5c28;
// ram_cell[     269] = 32'h0f0009c7;
// ram_cell[     270] = 32'hb5c4a293;
// ram_cell[     271] = 32'hb823ad8e;
// ram_cell[     272] = 32'h4d76a25d;
// ram_cell[     273] = 32'h30eb7e8d;
// ram_cell[     274] = 32'h3bb787f4;
// ram_cell[     275] = 32'he3b781fd;
// ram_cell[     276] = 32'h4b30362b;
// ram_cell[     277] = 32'h61059d1e;
// ram_cell[     278] = 32'h997bd92f;
// ram_cell[     279] = 32'h6fded37c;
// ram_cell[     280] = 32'hefc9dd8b;
// ram_cell[     281] = 32'h16389fea;
// ram_cell[     282] = 32'h9440997b;
// ram_cell[     283] = 32'h6a0b0f84;
// ram_cell[     284] = 32'h3bc2aa5e;
// ram_cell[     285] = 32'hd755a9d3;
// ram_cell[     286] = 32'h5343e57d;
// ram_cell[     287] = 32'he64da363;
// ram_cell[     288] = 32'h0b144b9a;
// ram_cell[     289] = 32'h4025e0ac;
// ram_cell[     290] = 32'h8955a025;
// ram_cell[     291] = 32'h4deaaec7;
// ram_cell[     292] = 32'he8f8c2ba;
// ram_cell[     293] = 32'h9e67db97;
// ram_cell[     294] = 32'h7ec3cef8;
// ram_cell[     295] = 32'he079b906;
// ram_cell[     296] = 32'h6d929e35;
// ram_cell[     297] = 32'he43971b4;
// ram_cell[     298] = 32'h09d5c098;
// ram_cell[     299] = 32'hf609e462;
// ram_cell[     300] = 32'hcff0fcd6;
// ram_cell[     301] = 32'h908cbaf3;
// ram_cell[     302] = 32'hb18c1185;
// ram_cell[     303] = 32'h1a46b9a9;
// ram_cell[     304] = 32'h4f8fdd8e;
// ram_cell[     305] = 32'h675a8e70;
// ram_cell[     306] = 32'h970bac6c;
// ram_cell[     307] = 32'hffe9b29e;
// ram_cell[     308] = 32'h92498fea;
// ram_cell[     309] = 32'h52ade204;
// ram_cell[     310] = 32'h3559918a;
// ram_cell[     311] = 32'h67fc367f;
// ram_cell[     312] = 32'hc423f655;
// ram_cell[     313] = 32'h0e1e964c;
// ram_cell[     314] = 32'h317e2c10;
// ram_cell[     315] = 32'h525986f0;
// ram_cell[     316] = 32'h38701a80;
// ram_cell[     317] = 32'h2354b798;
// ram_cell[     318] = 32'hd50e3dda;
// ram_cell[     319] = 32'hc4976532;
// ram_cell[     320] = 32'h0650de9f;
// ram_cell[     321] = 32'h65002110;
// ram_cell[     322] = 32'h5f4da4df;
// ram_cell[     323] = 32'h61d46659;
// ram_cell[     324] = 32'h19fe0d3b;
// ram_cell[     325] = 32'h0bfd0adc;
// ram_cell[     326] = 32'heda5c643;
// ram_cell[     327] = 32'hab07d154;
// ram_cell[     328] = 32'hb4379d17;
// ram_cell[     329] = 32'h8f63efe4;
// ram_cell[     330] = 32'hba981c2e;
// ram_cell[     331] = 32'h88708d28;
// ram_cell[     332] = 32'h28768765;
// ram_cell[     333] = 32'hb9cf248c;
// ram_cell[     334] = 32'hdcffdf2a;
// ram_cell[     335] = 32'hf10cb32b;
// ram_cell[     336] = 32'h6221abee;
// ram_cell[     337] = 32'hb2e66d77;
// ram_cell[     338] = 32'hfe2d68d5;
// ram_cell[     339] = 32'h635f526c;
// ram_cell[     340] = 32'h1aa24d71;
// ram_cell[     341] = 32'h4870cac8;
// ram_cell[     342] = 32'hcb650496;
// ram_cell[     343] = 32'h8ed01cf9;
// ram_cell[     344] = 32'he7936231;
// ram_cell[     345] = 32'hfbd30b25;
// ram_cell[     346] = 32'hc047cd0d;
// ram_cell[     347] = 32'h00685f8d;
// ram_cell[     348] = 32'h7cd480dc;
// ram_cell[     349] = 32'hd41d1456;
// ram_cell[     350] = 32'h6c9804b4;
// ram_cell[     351] = 32'hc6ff58e2;
// ram_cell[     352] = 32'h94da1ca4;
// ram_cell[     353] = 32'h9a60d05a;
// ram_cell[     354] = 32'h52bf51d8;
// ram_cell[     355] = 32'h61e4416f;
// ram_cell[     356] = 32'h2729f094;
// ram_cell[     357] = 32'hb3a8fdf8;
// ram_cell[     358] = 32'hb9a5f9d0;
// ram_cell[     359] = 32'hcabdb4f1;
// ram_cell[     360] = 32'h6410a604;
// ram_cell[     361] = 32'h7b2f7975;
// ram_cell[     362] = 32'h866444c9;
// ram_cell[     363] = 32'h3c405c46;
// ram_cell[     364] = 32'hbf6fe708;
// ram_cell[     365] = 32'hfba8911e;
// ram_cell[     366] = 32'h988f291d;
// ram_cell[     367] = 32'h633ab45f;
// ram_cell[     368] = 32'h93823e78;
// ram_cell[     369] = 32'h2211e650;
// ram_cell[     370] = 32'h669f10c8;
// ram_cell[     371] = 32'hba86df95;
// ram_cell[     372] = 32'h6fa932a0;
// ram_cell[     373] = 32'hfe198451;
// ram_cell[     374] = 32'h729ea642;
// ram_cell[     375] = 32'h1252b6db;
// ram_cell[     376] = 32'hba27c64d;
// ram_cell[     377] = 32'hbf4a4ff8;
// ram_cell[     378] = 32'h20eb45da;
// ram_cell[     379] = 32'h122023da;
// ram_cell[     380] = 32'h1b01b97b;
// ram_cell[     381] = 32'h44619ead;
// ram_cell[     382] = 32'h62cfb4fa;
// ram_cell[     383] = 32'hd8c12730;
// ram_cell[     384] = 32'ha6268cdc;
// ram_cell[     385] = 32'h00757d3a;
// ram_cell[     386] = 32'hd62f86e5;
// ram_cell[     387] = 32'hfe5ee57c;
// ram_cell[     388] = 32'h3179a2d6;
// ram_cell[     389] = 32'h2da6d88b;
// ram_cell[     390] = 32'hc1e73f0a;
// ram_cell[     391] = 32'h2b8e52d7;
// ram_cell[     392] = 32'h3a662409;
// ram_cell[     393] = 32'h8e701389;
// ram_cell[     394] = 32'h6d90351d;
// ram_cell[     395] = 32'h76243b15;
// ram_cell[     396] = 32'hff787dbf;
// ram_cell[     397] = 32'h442aa0a6;
// ram_cell[     398] = 32'hb5fc30be;
// ram_cell[     399] = 32'h9626ef22;
// ram_cell[     400] = 32'he1a8c6b4;
// ram_cell[     401] = 32'hd6f5ec70;
// ram_cell[     402] = 32'h157d9ffc;
// ram_cell[     403] = 32'h4c61c664;
// ram_cell[     404] = 32'hcf03646e;
// ram_cell[     405] = 32'h942c4ecd;
// ram_cell[     406] = 32'h119de4bd;
// ram_cell[     407] = 32'h6a5190b4;
// ram_cell[     408] = 32'h32cf8eba;
// ram_cell[     409] = 32'h20d6061a;
// ram_cell[     410] = 32'h6fffd9e3;
// ram_cell[     411] = 32'hd93f8dac;
// ram_cell[     412] = 32'h456f03ec;
// ram_cell[     413] = 32'hc8efdaf1;
// ram_cell[     414] = 32'h866eb62b;
// ram_cell[     415] = 32'h81dc2edd;
// ram_cell[     416] = 32'h5d2ab490;
// ram_cell[     417] = 32'h2584cf40;
// ram_cell[     418] = 32'h543b262f;
// ram_cell[     419] = 32'h7d75707b;
// ram_cell[     420] = 32'h08f95980;
// ram_cell[     421] = 32'hbd124b49;
// ram_cell[     422] = 32'hef504470;
// ram_cell[     423] = 32'hae5460d3;
// ram_cell[     424] = 32'h78cb0ba9;
// ram_cell[     425] = 32'hc300ff50;
// ram_cell[     426] = 32'he9ad99f6;
// ram_cell[     427] = 32'hb630768d;
// ram_cell[     428] = 32'hea7fdaed;
// ram_cell[     429] = 32'he48fa5f6;
// ram_cell[     430] = 32'h13a2812b;
// ram_cell[     431] = 32'h0b18aa88;
// ram_cell[     432] = 32'hc6ccd3c4;
// ram_cell[     433] = 32'hfc4f3856;
// ram_cell[     434] = 32'hd500b530;
// ram_cell[     435] = 32'h45fb1fde;
// ram_cell[     436] = 32'h6f86ea7f;
// ram_cell[     437] = 32'h666702dc;
// ram_cell[     438] = 32'hde994d5b;
// ram_cell[     439] = 32'h5815c634;
// ram_cell[     440] = 32'ha986cf04;
// ram_cell[     441] = 32'h442b9775;
// ram_cell[     442] = 32'he2d0ca1a;
// ram_cell[     443] = 32'h88ee0f4d;
// ram_cell[     444] = 32'h6aa8f69a;
// ram_cell[     445] = 32'h1bf8d023;
// ram_cell[     446] = 32'h8ee60e12;
// ram_cell[     447] = 32'h1f6a5891;
// ram_cell[     448] = 32'h4a2ca347;
// ram_cell[     449] = 32'h71e051ba;
// ram_cell[     450] = 32'hc67500f9;
// ram_cell[     451] = 32'h41ed9a85;
// ram_cell[     452] = 32'h5be7a7c4;
// ram_cell[     453] = 32'h2dd825d5;
// ram_cell[     454] = 32'h598abde9;
// ram_cell[     455] = 32'h447d1bbb;
// ram_cell[     456] = 32'h35edcb3c;
// ram_cell[     457] = 32'hb971d1e8;
// ram_cell[     458] = 32'h1f80fbea;
// ram_cell[     459] = 32'hcd617e98;
// ram_cell[     460] = 32'h0446c058;
// ram_cell[     461] = 32'h38e400f9;
// ram_cell[     462] = 32'h6ddd8f24;
// ram_cell[     463] = 32'h5b609feb;
// ram_cell[     464] = 32'h56c7271a;
// ram_cell[     465] = 32'h3eed45f2;
// ram_cell[     466] = 32'h729d9ce6;
// ram_cell[     467] = 32'h969e7eb9;
// ram_cell[     468] = 32'h9e0482b7;
// ram_cell[     469] = 32'h294a58c6;
// ram_cell[     470] = 32'h3b7f5794;
// ram_cell[     471] = 32'h7efc19cd;
// ram_cell[     472] = 32'hf4738a60;
// ram_cell[     473] = 32'he129effe;
// ram_cell[     474] = 32'h905beb88;
// ram_cell[     475] = 32'he3a3b93b;
// ram_cell[     476] = 32'hf6e4434e;
// ram_cell[     477] = 32'h030ce8ac;
// ram_cell[     478] = 32'h57133b1d;
// ram_cell[     479] = 32'h6926ff49;
// ram_cell[     480] = 32'hc71b38c2;
// ram_cell[     481] = 32'h4ff063f7;
// ram_cell[     482] = 32'h94cbe140;
// ram_cell[     483] = 32'hddf786da;
// ram_cell[     484] = 32'hde13539b;
// ram_cell[     485] = 32'h1bae2906;
// ram_cell[     486] = 32'h4989f21a;
// ram_cell[     487] = 32'h130a72ac;
// ram_cell[     488] = 32'h8772f34c;
// ram_cell[     489] = 32'h688a7154;
// ram_cell[     490] = 32'h71a75c66;
// ram_cell[     491] = 32'h68c0c449;
// ram_cell[     492] = 32'hd2ecfefb;
// ram_cell[     493] = 32'h8cf14fc1;
// ram_cell[     494] = 32'hf4290d9a;
// ram_cell[     495] = 32'h525a2758;
// ram_cell[     496] = 32'h7c1c8f7d;
// ram_cell[     497] = 32'hd09a14a5;
// ram_cell[     498] = 32'hb1ffc2c6;
// ram_cell[     499] = 32'hdc8e4969;
// ram_cell[     500] = 32'hb03d0347;
// ram_cell[     501] = 32'hb26afb7d;
// ram_cell[     502] = 32'h9db27864;
// ram_cell[     503] = 32'h41ee9331;
// ram_cell[     504] = 32'hc386058d;
// ram_cell[     505] = 32'hc2164ff3;
// ram_cell[     506] = 32'hfe18ae8d;
// ram_cell[     507] = 32'hea7fc8ee;
// ram_cell[     508] = 32'h031b2d6b;
// ram_cell[     509] = 32'h1dc30c0f;
// ram_cell[     510] = 32'hd3b94b6e;
// ram_cell[     511] = 32'h3cd2b778;
// // src matrix B
// ram_cell[     512] = 32'h5337fca8;
// ram_cell[     513] = 32'h8ac3642f;
// ram_cell[     514] = 32'hfd3a1f8f;
// ram_cell[     515] = 32'hc2f33a6f;
// ram_cell[     516] = 32'h7c68613d;
// ram_cell[     517] = 32'h9a2a7482;
// ram_cell[     518] = 32'ha145e3e6;
// ram_cell[     519] = 32'ha7a10a31;
// ram_cell[     520] = 32'h347bf859;
// ram_cell[     521] = 32'hc93938d4;
// ram_cell[     522] = 32'hed7d4cb8;
// ram_cell[     523] = 32'hee6d8cd2;
// ram_cell[     524] = 32'hfea6156c;
// ram_cell[     525] = 32'h0746e83b;
// ram_cell[     526] = 32'h68925033;
// ram_cell[     527] = 32'h8312a1b2;
// ram_cell[     528] = 32'h24f1dc36;
// ram_cell[     529] = 32'h1436952e;
// ram_cell[     530] = 32'hc2103b29;
// ram_cell[     531] = 32'h1cac9599;
// ram_cell[     532] = 32'h737b032d;
// ram_cell[     533] = 32'h64a8cf4c;
// ram_cell[     534] = 32'hfe2be210;
// ram_cell[     535] = 32'he0b96947;
// ram_cell[     536] = 32'hacb0aa21;
// ram_cell[     537] = 32'h3da6a64f;
// ram_cell[     538] = 32'h6ae2bf07;
// ram_cell[     539] = 32'h61d83fb7;
// ram_cell[     540] = 32'h3121ecda;
// ram_cell[     541] = 32'h40faf598;
// ram_cell[     542] = 32'hc2fd2713;
// ram_cell[     543] = 32'h8aa07bf4;
// ram_cell[     544] = 32'h97428230;
// ram_cell[     545] = 32'h758dfb96;
// ram_cell[     546] = 32'h0b42a890;
// ram_cell[     547] = 32'h1ed6ce15;
// ram_cell[     548] = 32'h9fff5900;
// ram_cell[     549] = 32'hd45ace77;
// ram_cell[     550] = 32'h2172f7cd;
// ram_cell[     551] = 32'hbcabc1a3;
// ram_cell[     552] = 32'he5f86e01;
// ram_cell[     553] = 32'hb7057b36;
// ram_cell[     554] = 32'hf55e1ffe;
// ram_cell[     555] = 32'h8075552b;
// ram_cell[     556] = 32'h3c56a995;
// ram_cell[     557] = 32'h16c7ff4d;
// ram_cell[     558] = 32'h7fe529bd;
// ram_cell[     559] = 32'h34ef1ba4;
// ram_cell[     560] = 32'hf4c6458a;
// ram_cell[     561] = 32'h43beeaf0;
// ram_cell[     562] = 32'h37ee97b7;
// ram_cell[     563] = 32'haf054ba1;
// ram_cell[     564] = 32'h62e5506d;
// ram_cell[     565] = 32'h38915b1a;
// ram_cell[     566] = 32'h391ecc67;
// ram_cell[     567] = 32'h568b7068;
// ram_cell[     568] = 32'h1b98267e;
// ram_cell[     569] = 32'hbab2f710;
// ram_cell[     570] = 32'hcb76e8dc;
// ram_cell[     571] = 32'ha3e84639;
// ram_cell[     572] = 32'h8bafc414;
// ram_cell[     573] = 32'h3f2bed8c;
// ram_cell[     574] = 32'h349d1118;
// ram_cell[     575] = 32'hc3829765;
// ram_cell[     576] = 32'h286f8d17;
// ram_cell[     577] = 32'hffbbc576;
// ram_cell[     578] = 32'hb3bad8dc;
// ram_cell[     579] = 32'hddccad57;
// ram_cell[     580] = 32'h7f993f2d;
// ram_cell[     581] = 32'h55c23787;
// ram_cell[     582] = 32'h99b6fb64;
// ram_cell[     583] = 32'h3dbba321;
// ram_cell[     584] = 32'hb2285104;
// ram_cell[     585] = 32'had13db26;
// ram_cell[     586] = 32'h736f2738;
// ram_cell[     587] = 32'hd33386dd;
// ram_cell[     588] = 32'h649f61d5;
// ram_cell[     589] = 32'ha4244adf;
// ram_cell[     590] = 32'ha859505b;
// ram_cell[     591] = 32'hee3f77b8;
// ram_cell[     592] = 32'ha91930e5;
// ram_cell[     593] = 32'h1e52b157;
// ram_cell[     594] = 32'h7c48a3c5;
// ram_cell[     595] = 32'h4701596e;
// ram_cell[     596] = 32'h1703fabe;
// ram_cell[     597] = 32'h469f6251;
// ram_cell[     598] = 32'hc7dd4490;
// ram_cell[     599] = 32'he517f92b;
// ram_cell[     600] = 32'h73549394;
// ram_cell[     601] = 32'hc7a802bd;
// ram_cell[     602] = 32'h0be954a0;
// ram_cell[     603] = 32'h205f5eee;
// ram_cell[     604] = 32'h55ed1079;
// ram_cell[     605] = 32'h30823162;
// ram_cell[     606] = 32'h7f0d9208;
// ram_cell[     607] = 32'hab163dfe;
// ram_cell[     608] = 32'h0f139081;
// ram_cell[     609] = 32'h5eeb6954;
// ram_cell[     610] = 32'hb23b015e;
// ram_cell[     611] = 32'h4e21c654;
// ram_cell[     612] = 32'hb74c28f9;
// ram_cell[     613] = 32'h88573170;
// ram_cell[     614] = 32'h09987ed3;
// ram_cell[     615] = 32'h863038fc;
// ram_cell[     616] = 32'hef102ee9;
// ram_cell[     617] = 32'ha5d4ad7c;
// ram_cell[     618] = 32'h4b974719;
// ram_cell[     619] = 32'h5ec921a1;
// ram_cell[     620] = 32'h6e5962cd;
// ram_cell[     621] = 32'h38bca434;
// ram_cell[     622] = 32'h373f2ecb;
// ram_cell[     623] = 32'h275bb394;
// ram_cell[     624] = 32'he9688334;
// ram_cell[     625] = 32'h0d688a68;
// ram_cell[     626] = 32'h29848b3e;
// ram_cell[     627] = 32'hfac9f56b;
// ram_cell[     628] = 32'h444db862;
// ram_cell[     629] = 32'hce7ab8e2;
// ram_cell[     630] = 32'h9524961c;
// ram_cell[     631] = 32'h64d5d665;
// ram_cell[     632] = 32'he9cf3b5b;
// ram_cell[     633] = 32'h64456148;
// ram_cell[     634] = 32'h7165a076;
// ram_cell[     635] = 32'h1ffc48cc;
// ram_cell[     636] = 32'ha2dd4cd5;
// ram_cell[     637] = 32'h1fff4dcb;
// ram_cell[     638] = 32'h2f6e2efd;
// ram_cell[     639] = 32'h26920a13;
// ram_cell[     640] = 32'ha547abba;
// ram_cell[     641] = 32'h9ab85120;
// ram_cell[     642] = 32'ha3e22ec1;
// ram_cell[     643] = 32'hf2969870;
// ram_cell[     644] = 32'h498f323a;
// ram_cell[     645] = 32'h890cb9e3;
// ram_cell[     646] = 32'h1fe602ce;
// ram_cell[     647] = 32'h120110cf;
// ram_cell[     648] = 32'h7b747eb3;
// ram_cell[     649] = 32'hfae36867;
// ram_cell[     650] = 32'hef6e64eb;
// ram_cell[     651] = 32'h8b54d5b5;
// ram_cell[     652] = 32'ha5dc94c2;
// ram_cell[     653] = 32'hf1185082;
// ram_cell[     654] = 32'h1505886e;
// ram_cell[     655] = 32'hd177885f;
// ram_cell[     656] = 32'he66539cc;
// ram_cell[     657] = 32'h2665e768;
// ram_cell[     658] = 32'h2958266a;
// ram_cell[     659] = 32'h1bc35b75;
// ram_cell[     660] = 32'h67ed4e93;
// ram_cell[     661] = 32'h0ba84e27;
// ram_cell[     662] = 32'hed14a8c6;
// ram_cell[     663] = 32'haf1b3df2;
// ram_cell[     664] = 32'h8f536108;
// ram_cell[     665] = 32'haf24a9c9;
// ram_cell[     666] = 32'h039e5638;
// ram_cell[     667] = 32'ha72d8c0b;
// ram_cell[     668] = 32'h0f19120b;
// ram_cell[     669] = 32'h835bc7f3;
// ram_cell[     670] = 32'h81f6b173;
// ram_cell[     671] = 32'hbc79f6fd;
// ram_cell[     672] = 32'h28400f39;
// ram_cell[     673] = 32'haff536df;
// ram_cell[     674] = 32'h080a34cb;
// ram_cell[     675] = 32'h6d977bde;
// ram_cell[     676] = 32'h12267b80;
// ram_cell[     677] = 32'h5235637d;
// ram_cell[     678] = 32'h589f217f;
// ram_cell[     679] = 32'h193c5ee9;
// ram_cell[     680] = 32'hd3ed127d;
// ram_cell[     681] = 32'h0b0d6a2f;
// ram_cell[     682] = 32'h4a9bdc7c;
// ram_cell[     683] = 32'hb1a833f1;
// ram_cell[     684] = 32'had4b999c;
// ram_cell[     685] = 32'h9ec9076e;
// ram_cell[     686] = 32'h2d3e4e22;
// ram_cell[     687] = 32'hb902a387;
// ram_cell[     688] = 32'he830ffee;
// ram_cell[     689] = 32'h9a7bf93d;
// ram_cell[     690] = 32'h0287726f;
// ram_cell[     691] = 32'h21b407f9;
// ram_cell[     692] = 32'h47d3ee57;
// ram_cell[     693] = 32'h782caf5c;
// ram_cell[     694] = 32'h7d42ece4;
// ram_cell[     695] = 32'hb2a06d28;
// ram_cell[     696] = 32'ha41f7f8e;
// ram_cell[     697] = 32'h63ac0cbe;
// ram_cell[     698] = 32'h87213209;
// ram_cell[     699] = 32'h7d950b0a;
// ram_cell[     700] = 32'h5df905f8;
// ram_cell[     701] = 32'hd50e0dac;
// ram_cell[     702] = 32'h85ac37fc;
// ram_cell[     703] = 32'hc00b8a2c;
// ram_cell[     704] = 32'h7372731d;
// ram_cell[     705] = 32'h22b1b6ee;
// ram_cell[     706] = 32'hfb08f9be;
// ram_cell[     707] = 32'h1c242e94;
// ram_cell[     708] = 32'h08b85e74;
// ram_cell[     709] = 32'h0e899c57;
// ram_cell[     710] = 32'h5e46c081;
// ram_cell[     711] = 32'h5b7d4776;
// ram_cell[     712] = 32'he40090ff;
// ram_cell[     713] = 32'h6b5e117c;
// ram_cell[     714] = 32'h7d8baba0;
// ram_cell[     715] = 32'hd5567f16;
// ram_cell[     716] = 32'h2a839f67;
// ram_cell[     717] = 32'hc3ca8e11;
// ram_cell[     718] = 32'he92f48c5;
// ram_cell[     719] = 32'h8479f843;
// ram_cell[     720] = 32'h50c05ee5;
// ram_cell[     721] = 32'h48b63cfa;
// ram_cell[     722] = 32'h7cd8ff20;
// ram_cell[     723] = 32'hb60ad992;
// ram_cell[     724] = 32'h1e8b48ef;
// ram_cell[     725] = 32'hfa57a284;
// ram_cell[     726] = 32'h75b7ee53;
// ram_cell[     727] = 32'h8e847b8a;
// ram_cell[     728] = 32'hd2a584f9;
// ram_cell[     729] = 32'h20811860;
// ram_cell[     730] = 32'h7619db3b;
// ram_cell[     731] = 32'h102fea52;
// ram_cell[     732] = 32'h215dd570;
// ram_cell[     733] = 32'h8c29a689;
// ram_cell[     734] = 32'h17fad848;
// ram_cell[     735] = 32'h5c9073b8;
// ram_cell[     736] = 32'h0b833e89;
// ram_cell[     737] = 32'h3ff3ba21;
// ram_cell[     738] = 32'h39bee887;
// ram_cell[     739] = 32'h02fecefa;
// ram_cell[     740] = 32'h73fb8112;
// ram_cell[     741] = 32'h95c82a46;
// ram_cell[     742] = 32'hd0c9bdaf;
// ram_cell[     743] = 32'hf74b89e2;
// ram_cell[     744] = 32'ha3affa77;
// ram_cell[     745] = 32'h3286c6f8;
// ram_cell[     746] = 32'h26c8b346;
// ram_cell[     747] = 32'h45754d8b;
// ram_cell[     748] = 32'h1d9169d0;
// ram_cell[     749] = 32'h0f2332be;
// ram_cell[     750] = 32'h016ba687;
// ram_cell[     751] = 32'h7c9e3800;
// ram_cell[     752] = 32'hf4eff073;
// ram_cell[     753] = 32'h902254d7;
// ram_cell[     754] = 32'h9aa5a923;
// ram_cell[     755] = 32'hd28d03be;
// ram_cell[     756] = 32'h5a85791b;
// ram_cell[     757] = 32'h102c83f5;
// ram_cell[     758] = 32'h8e7c8503;
// ram_cell[     759] = 32'h07248bab;
// ram_cell[     760] = 32'hbde4754e;
// ram_cell[     761] = 32'he8c3ee57;
// ram_cell[     762] = 32'h7cafc551;
// ram_cell[     763] = 32'h1c89d67b;
// ram_cell[     764] = 32'h817158c1;
// ram_cell[     765] = 32'hdf4f757f;
// ram_cell[     766] = 32'head1a369;
// ram_cell[     767] = 32'h17e149c7;
// end

// endmodule



