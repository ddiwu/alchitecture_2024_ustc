�� 
 m o d u l e   m e m   # (                                       / /    
         p a r a m e t e r     A D D R _ L E N     =   1 1       / /    
 )   (  
         i n p u t     c l k ,   r s t ,  
         i n p u t     [ A D D R _ L E N - 1 : 0 ]   a d d r ,   / /   m e m o r y   a d d r e s s  
         o u t p u t   r e g   [ 3 1 : 0 ]   r d _ d a t a ,     / /   d a t a   r e a d   o u t  
         i n p u t     w r _ r e q ,  
         i n p u t     [ 3 1 : 0 ]   w r _ d a t a               / /   d a t a   w r i t e   i n  
 ) ;  
 l o c a l p a r a m   M E M _ S I Z E   =   1 < < A D D R _ L E N ;  
 r e g   [ 3 1 : 0 ]   r a m _ c e l l   [ M E M _ S I Z E ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )  
                 r d _ d a t a   < =   0 ;  
         e l s e  
                 r d _ d a t a   < =   r a m _ c e l l [ a d d r ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k )  
         i f ( w r _ r e q )    
                 r a m _ c e l l [ a d d r ]   < =   w r _ d a t a ;  
  
 i n i t i a l   b e g i n  
         r a m _ c e l l [               0 ]   =   3 2 ' h 0 0 0 0 0 0 3 7 ;  
         r a m _ c e l l [               1 ]   =   3 2 ' h 0 0 0 0 0 0 a 6 ;  
         r a m _ c e l l [               2 ]   =   3 2 ' h 0 0 0 0 0 1 0 6 ;  
         r a m _ c e l l [               3 ]   =   3 2 ' h 0 0 0 0 0 0 7 0 ;  
         r a m _ c e l l [               4 ]   =   3 2 ' h 0 0 0 0 0 1 8 2 ;  
         r a m _ c e l l [               5 ]   =   3 2 ' h 0 0 0 0 0 1 7 8 ;  
         r a m _ c e l l [               6 ]   =   3 2 ' h 0 0 0 0 0 1 9 1 ;  
         r a m _ c e l l [               7 ]   =   3 2 ' h 0 0 0 0 0 0 9 f ;  
         r a m _ c e l l [               8 ]   =   3 2 ' h 0 0 0 0 0 1 e 6 ;  
         r a m _ c e l l [               9 ]   =   3 2 ' h 0 0 0 0 0 0 f 6 ;  
         r a m _ c e l l [             1 0 ]   =   3 2 ' h 0 0 0 0 0 1 2 f ;  
         r a m _ c e l l [             1 1 ]   =   3 2 ' h 0 0 0 0 0 1 4 3 ;  
         r a m _ c e l l [             1 2 ]   =   3 2 ' h 0 0 0 0 0 0 b 0 ;  
         r a m _ c e l l [             1 3 ]   =   3 2 ' h 0 0 0 0 0 1 1 4 ;  
         r a m _ c e l l [             1 4 ]   =   3 2 ' h 0 0 0 0 0 1 0 2 ;  
         r a m _ c e l l [             1 5 ]   =   3 2 ' h 0 0 0 0 0 0 b a ;  
         r a m _ c e l l [             1 6 ]   =   3 2 ' h 0 0 0 0 0 1 a 6 ;  
         r a m _ c e l l [             1 7 ]   =   3 2 ' h 0 0 0 0 0 0 b 3 ;  
         r a m _ c e l l [             1 8 ]   =   3 2 ' h 0 0 0 0 0 0 0 6 ;  
         r a m _ c e l l [             1 9 ]   =   3 2 ' h 0 0 0 0 0 0 7 9 ;  
         r a m _ c e l l [             2 0 ]   =   3 2 ' h 0 0 0 0 0 0 3 2 ;  
         r a m _ c e l l [             2 1 ]   =   3 2 ' h 0 0 0 0 0 1 d 0 ;  
         r a m _ c e l l [             2 2 ]   =   3 2 ' h 0 0 0 0 0 0 e 6 ;  
         r a m _ c e l l [             2 3 ]   =   3 2 ' h 0 0 0 0 0 0 0 1 ;  
         r a m _ c e l l [             2 4 ]   =   3 2 ' h 0 0 0 0 0 1 e 2 ;  
         r a m _ c e l l [             2 5 ]   =   3 2 ' h 0 0 0 0 0 1 f 3 ;  
         r a m _ c e l l [             2 6 ]   =   3 2 ' h 0 0 0 0 0 1 2 8 ;  
         r a m _ c e l l [             2 7 ]   =   3 2 ' h 0 0 0 0 0 0 9 e ;  
         r a m _ c e l l [             2 8 ]   =   3 2 ' h 0 0 0 0 0 1 0 b ;  
         r a m _ c e l l [             2 9 ]   =   3 2 ' h 0 0 0 0 0 1 b f ;  
         r a m _ c e l l [             3 0 ]   =   3 2 ' h 0 0 0 0 0 0 b 8 ;  
         r a m _ c e l l [             3 1 ]   =   3 2 ' h 0 0 0 0 0 1 4 0 ;  
         r a m _ c e l l [             3 2 ]   =   3 2 ' h 0 0 0 0 0 0 f d ;  
         r a m _ c e l l [             3 3 ]   =   3 2 ' h 0 0 0 0 0 1 f 9 ;  
         r a m _ c e l l [             3 4 ]   =   3 2 ' h 0 0 0 0 0 1 a d ;  
         r a m _ c e l l [             3 5 ]   =   3 2 ' h 0 0 0 0 0 0 0 3 ;  
         r a m _ c e l l [             3 6 ]   =   3 2 ' h 0 0 0 0 0 0 e 5 ;  
         r a m _ c e l l [             3 7 ]   =   3 2 ' h 0 0 0 0 0 1 f 2 ;  
         r a m _ c e l l [             3 8 ]   =   3 2 ' h 0 0 0 0 0 1 d 9 ;  
         r a m _ c e l l [             3 9 ]   =   3 2 ' h 0 0 0 0 0 0 f b ;  
         r a m _ c e l l [             4 0 ]   =   3 2 ' h 0 0 0 0 0 1 9 9 ;  
         r a m _ c e l l [             4 1 ]   =   3 2 ' h 0 0 0 0 0 1 e 8 ;  
         r a m _ c e l l [             4 2 ]   =   3 2 ' h 0 0 0 0 0 0 2 9 ;  
         r a m _ c e l l [             4 3 ]   =   3 2 ' h 0 0 0 0 0 1 7 9 ;  
         r a m _ c e l l [             4 4 ]   =   3 2 ' h 0 0 0 0 0 0 4 8 ;  
         r a m _ c e l l [             4 5 ]   =   3 2 ' h 0 0 0 0 0 0 a b ;  
         r a m _ c e l l [             4 6 ]   =   3 2 ' h 0 0 0 0 0 0 c a ;  
         r a m _ c e l l [             4 7 ]   =   3 2 ' h 0 0 0 0 0 0 9 2 ;  
         r a m _ c e l l [             4 8 ]   =   3 2 ' h 0 0 0 0 0 1 b 3 ;  
         r a m _ c e l l [             4 9 ]   =   3 2 ' h 0 0 0 0 0 0 a 8 ;  
         r a m _ c e l l [             5 0 ]   =   3 2 ' h 0 0 0 0 0 1 b 9 ;  
         r a m _ c e l l [             5 1 ]   =   3 2 ' h 0 0 0 0 0 1 f 6 ;  
         r a m _ c e l l [             5 2 ]   =   3 2 ' h 0 0 0 0 0 1 d b ;  
         r a m _ c e l l [             5 3 ]   =   3 2 ' h 0 0 0 0 0 0 8 7 ;  
         r a m _ c e l l [             5 4 ]   =   3 2 ' h 0 0 0 0 0 1 6 3 ;  
         r a m _ c e l l [             5 5 ]   =   3 2 ' h 0 0 0 0 0 1 b 0 ;  
         r a m _ c e l l [             5 6 ]   =   3 2 ' h 0 0 0 0 0 1 8 5 ;  
         r a m _ c e l l [             5 7 ]   =   3 2 ' h 0 0 0 0 0 1 a f ;  
         r a m _ c e l l [             5 8 ]   =   3 2 ' h 0 0 0 0 0 1 c 9 ;  
         r a m _ c e l l [             5 9 ]   =   3 2 ' h 0 0 0 0 0 1 4 8 ;  
         r a m _ c e l l [             6 0 ]   =   3 2 ' h 0 0 0 0 0 1 8 f ;  
         r a m _ c e l l [             6 1 ]   =   3 2 ' h 0 0 0 0 0 1 8 6 ;  
         r a m _ c e l l [             6 2 ]   =   3 2 ' h 0 0 0 0 0 0 1 f ;  
         r a m _ c e l l [             6 3 ]   =   3 2 ' h 0 0 0 0 0 0 3 c ;  
         r a m _ c e l l [             6 4 ]   =   3 2 ' h 0 0 0 0 0 1 4 2 ;  
         r a m _ c e l l [             6 5 ]   =   3 2 ' h 0 0 0 0 0 1 6 4 ;  
         r a m _ c e l l [             6 6 ]   =   3 2 ' h 0 0 0 0 0 1 4 e ;  
         r a m _ c e l l [             6 7 ]   =   3 2 ' h 0 0 0 0 0 0 a f ;  
         r a m _ c e l l [             6 8 ]   =   3 2 ' h 0 0 0 0 0 0 9 7 ;  
         r a m _ c e l l [             6 9 ]   =   3 2 ' h 0 0 0 0 0 1 c 0 ;  
         r a m _ c e l l [             7 0 ]   =   3 2 ' h 0 0 0 0 0 1 7 f ;  
         r a m _ c e l l [             7 1 ]   =   3 2 ' h 0 0 0 0 0 1 7 5 ;  
         r a m _ c e l l [             7 2 ]   =   3 2 ' h 0 0 0 0 0 1 6 5 ;  
         r a m _ c e l l [             7 3 ]   =   3 2 ' h 0 0 0 0 0 1 3 8 ;  
         r a m _ c e l l [             7 4 ]   =   3 2 ' h 0 0 0 0 0 1 d e ;  
         r a m _ c e l l [             7 5 ]   =   3 2 ' h 0 0 0 0 0 0 0 c ;  
         r a m _ c e l l [             7 6 ]   =   3 2 ' h 0 0 0 0 0 0 6 5 ;  
         r a m _ c e l l [             7 7 ]   =   3 2 ' h 0 0 0 0 0 0 8 5 ;  
         r a m _ c e l l [             7 8 ]   =   3 2 ' h 0 0 0 0 0 0 3 1 ;  
         r a m _ c e l l [             7 9 ]   =   3 2 ' h 0 0 0 0 0 1 6 d ;  
         r a m _ c e l l [             8 0 ]   =   3 2 ' h 0 0 0 0 0 0 1 2 ;  
         r a m _ c e l l [             8 1 ]   =   3 2 ' h 0 0 0 0 0 0 4 a ;  
         r a m _ c e l l [             8 2 ]   =   3 2 ' h 0 0 0 0 0 0 5 5 ;  
         r a m _ c e l l [             8 3 ]   =   3 2 ' h 0 0 0 0 0 0 f 7 ;  
         r a m _ c e l l [             8 4 ]   =   3 2 ' h 0 0 0 0 0 1 4 1 ;  
         r a m _ c e l l [             8 5 ]   =   3 2 ' h 0 0 0 0 0 1 0 7 ;  
         r a m _ c e l l [             8 6 ]   =   3 2 ' h 0 0 0 0 0 1 1 2 ;  
         r a m _ c e l l [             8 7 ]   =   3 2 ' h 0 0 0 0 0 1 f 5 ;  
         r a m _ c e l l [             8 8 ]   =   3 2 ' h 0 0 0 0 0 1 d 1 ;  
         r a m _ c e l l [             8 9 ]   =   3 2 ' h 0 0 0 0 0 0 6 f ;  
         r a m _ c e l l [             9 0 ]   =   3 2 ' h 0 0 0 0 0 1 6 a ;  
         r a m _ c e l l [             9 1 ]   =   3 2 ' h 0 0 0 0 0 0 d b ;  
         r a m _ c e l l [             9 2 ]   =   3 2 ' h 0 0 0 0 0 1 5 c ;  
         r a m _ c e l l [             9 3 ]   =   3 2 ' h 0 0 0 0 0 0 0 b ;  
         r a m _ c e l l [             9 4 ]   =   3 2 ' h 0 0 0 0 0 1 c a ;  
         r a m _ c e l l [             9 5 ]   =   3 2 ' h 0 0 0 0 0 0 6 2 ;  
         r a m _ c e l l [             9 6 ]   =   3 2 ' h 0 0 0 0 0 1 5 9 ;  
         r a m _ c e l l [             9 7 ]   =   3 2 ' h 0 0 0 0 0 1 9 7 ;  
         r a m _ c e l l [             9 8 ]   =   3 2 ' h 0 0 0 0 0 1 5 f ;  
         r a m _ c e l l [             9 9 ]   =   3 2 ' h 0 0 0 0 0 1 b 4 ;  
         r a m _ c e l l [           1 0 0 ]   =   3 2 ' h 0 0 0 0 0 0 9 3 ;  
         r a m _ c e l l [           1 0 1 ]   =   3 2 ' h 0 0 0 0 0 1 e 9 ;  
         r a m _ c e l l [           1 0 2 ]   =   3 2 ' h 0 0 0 0 0 0 a 9 ;  
         r a m _ c e l l [           1 0 3 ]   =   3 2 ' h 0 0 0 0 0 1 1 1 ;  
         r a m _ c e l l [           1 0 4 ]   =   3 2 ' h 0 0 0 0 0 1 a 8 ;  
         r a m _ c e l l [           1 0 5 ]   =   3 2 ' h 0 0 0 0 0 0 f a ;  
         r a m _ c e l l [           1 0 6 ]   =   3 2 ' h 0 0 0 0 0 0 4 e ;  
         r a m _ c e l l [           1 0 7 ]   =   3 2 ' h 0 0 0 0 0 0 b 6 ;  
         r a m _ c e l l [           1 0 8 ]   =   3 2 ' h 0 0 0 0 0 0 c 2 ;  
         r a m _ c e l l [           1 0 9 ]   =   3 2 ' h 0 0 0 0 0 1 e d ;  
         r a m _ c e l l [           1 1 0 ]   =   3 2 ' h 0 0 0 0 0 0 0 e ;  
         r a m _ c e l l [           1 1 1 ]   =   3 2 ' h 0 0 0 0 0 1 0 3 ;  
         r a m _ c e l l [           1 1 2 ]   =   3 2 ' h 0 0 0 0 0 0 8 2 ;  
         r a m _ c e l l [           1 1 3 ]   =   3 2 ' h 0 0 0 0 0 1 6 2 ;  
         r a m _ c e l l [           1 1 4 ]   =   3 2 ' h 0 0 0 0 0 0 c e ;  
         r a m _ c e l l [           1 1 5 ]   =   3 2 ' h 0 0 0 0 0 1 2 4 ;  
         r a m _ c e l l [           1 1 6 ]   =   3 2 ' h 0 0 0 0 0 1 1 5 ;  
         r a m _ c e l l [           1 1 7 ]   =   3 2 ' h 0 0 0 0 0 0 d f ;  
         r a m _ c e l l [           1 1 8 ]   =   3 2 ' h 0 0 0 0 0 0 e 3 ;  
         r a m _ c e l l [           1 1 9 ]   =   3 2 ' h 0 0 0 0 0 1 2 e ;  
         r a m _ c e l l [           1 2 0 ]   =   3 2 ' h 0 0 0 0 0 1 c 3 ;  
         r a m _ c e l l [           1 2 1 ]   =   3 2 ' h 0 0 0 0 0 1 c 7 ;  
         r a m _ c e l l [           1 2 2 ]   =   3 2 ' h 0 0 0 0 0 1 a c ;  
         r a m _ c e l l [           1 2 3 ]   =   3 2 ' h 0 0 0 0 0 0 2 6 ;  
         r a m _ c e l l [           1 2 4 ]   =   3 2 ' h 0 0 0 0 0 0 4 c ;  
         r a m _ c e l l [           1 2 5 ]   =   3 2 ' h 0 0 0 0 0 1 0 8 ;  
         r a m _ c e l l [           1 2 6 ]   =   3 2 ' h 0 0 0 0 0 0 6 0 ;  
         r a m _ c e l l [           1 2 7 ]   =   3 2 ' h 0 0 0 0 0 0 b b ;  
         r a m _ c e l l [           1 2 8 ]   =   3 2 ' h 0 0 0 0 0 0 9 c ;  
         r a m _ c e l l [           1 2 9 ]   =   3 2 ' h 0 0 0 0 0 0 6 8 ;  
         r a m _ c e l l [           1 3 0 ]   =   3 2 ' h 0 0 0 0 0 0 3 3 ;  
         r a m _ c e l l [           1 3 1 ]   =   3 2 ' h 0 0 0 0 0 1 5 e ;  
         r a m _ c e l l [           1 3 2 ]   =   3 2 ' h 0 0 0 0 0 0 f 5 ;  
         r a m _ c e l l [           1 3 3 ]   =   3 2 ' h 0 0 0 0 0 1 9 5 ;  
         r a m _ c e l l [           1 3 4 ]   =   3 2 ' h 0 0 0 0 0 0 2 5 ;  
         r a m _ c e l l [           1 3 5 ]   =   3 2 ' h 0 0 0 0 0 0 1 8 ;  
         r a m _ c e l l [           1 3 6 ]   =   3 2 ' h 0 0 0 0 0 0 6 b ;  
         r a m _ c e l l [           1 3 7 ]   =   3 2 ' h 0 0 0 0 0 1 a 5 ;  
         r a m _ c e l l [           1 3 8 ]   =   3 2 ' h 0 0 0 0 0 1 4 7 ;  
         r a m _ c e l l [           1 3 9 ]   =   3 2 ' h 0 0 0 0 0 1 8 9 ;  
         r a m _ c e l l [           1 4 0 ]   =   3 2 ' h 0 0 0 0 0 1 3 2 ;  
         r a m _ c e l l [           1 4 1 ]   =   3 2 ' h 0 0 0 0 0 0 2 7 ;  
         r a m _ c e l l [           1 4 2 ]   =   3 2 ' h 0 0 0 0 0 1 3 5 ;  
         r a m _ c e l l [           1 4 3 ]   =   3 2 ' h 0 0 0 0 0 1 9 d ;  
         r a m _ c e l l [           1 4 4 ]   =   3 2 ' h 0 0 0 0 0 1 0 a ;  
         r a m _ c e l l [           1 4 5 ]   =   3 2 ' h 0 0 0 0 0 0 e e ;  
         r a m _ c e l l [           1 4 6 ]   =   3 2 ' h 0 0 0 0 0 1 6 b ;  
         r a m _ c e l l [           1 4 7 ]   =   3 2 ' h 0 0 0 0 0 1 5 8 ;  
         r a m _ c e l l [           1 4 8 ]   =   3 2 ' h 0 0 0 0 0 1 f 8 ;  
         r a m _ c e l l [           1 4 9 ]   =   3 2 ' h 0 0 0 0 0 1 0 9 ;  
         r a m _ c e l l [           1 5 0 ]   =   3 2 ' h 0 0 0 0 0 0 4 2 ;  
         r a m _ c e l l [           1 5 1 ]   =   3 2 ' h 0 0 0 0 0 0 2 e ;  
         r a m _ c e l l [           1 5 2 ]   =   3 2 ' h 0 0 0 0 0 0 8 3 ;  
         r a m _ c e l l [           1 5 3 ]   =   3 2 ' h 0 0 0 0 0 0 2 0 ;  
         r a m _ c e l l [           1 5 4 ]   =   3 2 ' h 0 0 0 0 0 1 b b ;  
         r a m _ c e l l [           1 5 5 ]   =   3 2 ' h 0 0 0 0 0 0 a 4 ;  
         r a m _ c e l l [           1 5 6 ]   =   3 2 ' h 0 0 0 0 0 1 e 3 ;  
         r a m _ c e l l [           1 5 7 ]   =   3 2 ' h 0 0 0 0 0 0 1 c ;  
         r a m _ c e l l [           1 5 8 ]   =   3 2 ' h 0 0 0 0 0 0 4 b ;  
         r a m _ c e l l [           1 5 9 ]   =   3 2 ' h 0 0 0 0 0 1 6 6 ;  
         r a m _ c e l l [           1 6 0 ]   =   3 2 ' h 0 0 0 0 0 0 5 6 ;  
         r a m _ c e l l [           1 6 1 ]   =   3 2 ' h 0 0 0 0 0 1 3 6 ;  
         r a m _ c e l l [           1 6 2 ]   =   3 2 ' h 0 0 0 0 0 0 5 c ;  
         r a m _ c e l l [           1 6 3 ]   =   3 2 ' h 0 0 0 0 0 0 6 7 ;  
         r a m _ c e l l [           1 6 4 ]   =   3 2 ' h 0 0 0 0 0 1 7 0 ;  
         r a m _ c e l l [           1 6 5 ]   =   3 2 ' h 0 0 0 0 0 0 e b ;  
         r a m _ c e l l [           1 6 6 ]   =   3 2 ' h 0 0 0 0 0 0 d 1 ;  
         r a m _ c e l l [           1 6 7 ]   =   3 2 ' h 0 0 0 0 0 0 1 4 ;  
         r a m _ c e l l [           1 6 8 ]   =   3 2 ' h 0 0 0 0 0 1 9 e ;  
         r a m _ c e l l [           1 6 9 ]   =   3 2 ' h 0 0 0 0 0 1 2 a ;  
         r a m _ c e l l [           1 7 0 ]   =   3 2 ' h 0 0 0 0 0 1 a e ;  
         r a m _ c e l l [           1 7 1 ]   =   3 2 ' h 0 0 0 0 0 1 5 6 ;  
         r a m _ c e l l [           1 7 2 ]   =   3 2 ' h 0 0 0 0 0 1 8 c ;  
         r a m _ c e l l [           1 7 3 ]   =   3 2 ' h 0 0 0 0 0 1 5 5 ;  
         r a m _ c e l l [           1 7 4 ]   =   3 2 ' h 0 0 0 0 0 1 1 a ;  
         r a m _ c e l l [           1 7 5 ]   =   3 2 ' h 0 0 0 0 0 1 4 d ;  
         r a m _ c e l l [           1 7 6 ]   =   3 2 ' h 0 0 0 0 0 0 b 9 ;  
         r a m _ c e l l [           1 7 7 ]   =   3 2 ' h 0 0 0 0 0 1 9 3 ;  
         r a m _ c e l l [           1 7 8 ]   =   3 2 ' h 0 0 0 0 0 0 0 d ;  
         r a m _ c e l l [           1 7 9 ]   =   3 2 ' h 0 0 0 0 0 1 c d ;  
         r a m _ c e l l [           1 8 0 ]   =   3 2 ' h 0 0 0 0 0 1 5 4 ;  
         r a m _ c e l l [           1 8 1 ]   =   3 2 ' h 0 0 0 0 0 0 d 5 ;  
         r a m _ c e l l [           1 8 2 ]   =   3 2 ' h 0 0 0 0 0 1 b 2 ;  
         r a m _ c e l l [           1 8 3 ]   =   3 2 ' h 0 0 0 0 0 0 4 4 ;  
         r a m _ c e l l [           1 8 4 ]   =   3 2 ' h 0 0 0 0 0 0 7 8 ;  
         r a m _ c e l l [           1 8 5 ]   =   3 2 ' h 0 0 0 0 0 0 6 1 ;  
         r a m _ c e l l [           1 8 6 ]   =   3 2 ' h 0 0 0 0 0 0 5 0 ;  
         r a m _ c e l l [           1 8 7 ]   =   3 2 ' h 0 0 0 0 0 0 5 4 ;  
         r a m _ c e l l [           1 8 8 ]   =   3 2 ' h 0 0 0 0 0 1 e 7 ;  
         r a m _ c e l l [           1 8 9 ]   =   3 2 ' h 0 0 0 0 0 0 5 e ;  
         r a m _ c e l l [           1 9 0 ]   =   3 2 ' h 0 0 0 0 0 1 8 a ;  
         r a m _ c e l l [           1 9 1 ]   =   3 2 ' h 0 0 0 0 0 1 2 1 ;  
         r a m _ c e l l [           1 9 2 ]   =   3 2 ' h 0 0 0 0 0 0 7 5 ;  
         r a m _ c e l l [           1 9 3 ]   =   3 2 ' h 0 0 0 0 0 0 c 5 ;  
         r a m _ c e l l [           1 9 4 ]   =   3 2 ' h 0 0 0 0 0 0 8 d ;  
         r a m _ c e l l [           1 9 5 ]   =   3 2 ' h 0 0 0 0 0 0 e a ;  
         r a m _ c e l l [           1 9 6 ]   =   3 2 ' h 0 0 0 0 0 1 8 0 ;  
         r a m _ c e l l [           1 9 7 ]   =   3 2 ' h 0 0 0 0 0 0 b 7 ;  
         r a m _ c e l l [           1 9 8 ]   =   3 2 ' h 0 0 0 0 0 0 d 7 ;  
         r a m _ c e l l [           1 9 9 ]   =   3 2 ' h 0 0 0 0 0 0 2 c ;  
         r a m _ c e l l [           2 0 0 ]   =   3 2 ' h 0 0 0 0 0 0 a e ;  
         r a m _ c e l l [           2 0 1 ]   =   3 2 ' h 0 0 0 0 0 1 c 1 ;  
         r a m _ c e l l [           2 0 2 ]   =   3 2 ' h 0 0 0 0 0 0 e d ;  
         r a m _ c e l l [           2 0 3 ]   =   3 2 ' h 0 0 0 0 0 1 8 e ;  
         r a m _ c e l l [           2 0 4 ]   =   3 2 ' h 0 0 0 0 0 1 1 8 ;  
         r a m _ c e l l [           2 0 5 ]   =   3 2 ' h 0 0 0 0 0 1 e 5 ;  
         r a m _ c e l l [           2 0 6 ]   =   3 2 ' h 0 0 0 0 0 1 e a ;  
         r a m _ c e l l [           2 0 7 ]   =   3 2 ' h 0 0 0 0 0 0 1 1 ;  
         r a m _ c e l l [           2 0 8 ]   =   3 2 ' h 0 0 0 0 0 1 d 2 ;  
         r a m _ c e l l [           2 0 9 ]   =   3 2 ' h 0 0 0 0 0 1 1 9 ;  
         r a m _ c e l l [           2 1 0 ]   =   3 2 ' h 0 0 0 0 0 1 5 d ;  
         r a m _ c e l l [           2 1 1 ]   =   3 2 ' h 0 0 0 0 0 1 1 3 ;  
         r a m _ c e l l [           2 1 2 ]   =   3 2 ' h 0 0 0 0 0 0 5 9 ;  
         r a m _ c e l l [           2 1 3 ]   =   3 2 ' h 0 0 0 0 0 0 c c ;  
         r a m _ c e l l [           2 1 4 ]   =   3 2 ' h 0 0 0 0 0 0 d 4 ;  
         r a m _ c e l l [           2 1 5 ]   =   3 2 ' h 0 0 0 0 0 1 1 0 ;  
         r a m _ c e l l [           2 1 6 ]   =   3 2 ' h 0 0 0 0 0 0 1 5 ;  
         r a m _ c e l l [           2 1 7 ]   =   3 2 ' h 0 0 0 0 0 0 e c ;  
         r a m _ c e l l [           2 1 8 ]   =   3 2 ' h 0 0 0 0 0 1 2 2 ;  
         r a m _ c e l l [           2 1 9 ]   =   3 2 ' h 0 0 0 0 0 0 5 1 ;  
         r a m _ c e l l [           2 2 0 ]   =   3 2 ' h 0 0 0 0 0 1 a a ;  
         r a m _ c e l l [           2 2 1 ]   =   3 2 ' h 0 0 0 0 0 1 2 0 ;  
         r a m _ c e l l [           2 2 2 ]   =   3 2 ' h 0 0 0 0 0 0 7 2 ;  
         r a m _ c e l l [           2 2 3 ]   =   3 2 ' h 0 0 0 0 0 1 e f ;  
         r a m _ c e l l [           2 2 4 ]   =   3 2 ' h 0 0 0 0 0 0 8 1 ;  
         r a m _ c e l l [           2 2 5 ]   =   3 2 ' h 0 0 0 0 0 0 f 9 ;  
         r a m _ c e l l [           2 2 6 ]   =   3 2 ' h 0 0 0 0 0 1 4 f ;  
         r a m _ c e l l [           2 2 7 ]   =   3 2 ' h 0 0 0 0 0 1 f c ;  
         r a m _ c e l l [           2 2 8 ]   =   3 2 ' h 0 0 0 0 0 0 c 7 ;  
         r a m _ c e l l [           2 2 9 ]   =   3 2 ' h 0 0 0 0 0 0 6 c ;  
         r a m _ c e l l [           2 3 0 ]   =   3 2 ' h 0 0 0 0 0 0 7 a ;  
         r a m _ c e l l [           2 3 1 ]   =   3 2 ' h 0 0 0 0 0 0 9 b ;  
         r a m _ c e l l [           2 3 2 ]   =   3 2 ' h 0 0 0 0 0 1 9 a ;  
         r a m _ c e l l [           2 3 3 ]   =   3 2 ' h 0 0 0 0 0 0 4 7 ;  
         r a m _ c e l l [           2 3 4 ]   =   3 2 ' h 0 0 0 0 0 1 e 0 ;  
         r a m _ c e l l [           2 3 5 ]   =   3 2 ' h 0 0 0 0 0 1 3 7 ;  
         r a m _ c e l l [           2 3 6 ]   =   3 2 ' h 0 0 0 0 0 0 0 4 ;  
         r a m _ c e l l [           2 3 7 ]   =   3 2 ' h 0 0 0 0 0 0 2 f ;  
         r a m _ c e l l [           2 3 8 ]   =   3 2 ' h 0 0 0 0 0 1 6 f ;  
         r a m _ c e l l [           2 3 9 ]   =   3 2 ' h 0 0 0 0 0 0 b d ;  
         r a m _ c e l l [           2 4 0 ]   =   3 2 ' h 0 0 0 0 0 0 3 5 ;  
         r a m _ c e l l [           2 4 1 ]   =   3 2 ' h 0 0 0 0 0 1 d f ;  
         r a m _ c e l l [           2 4 2 ]   =   3 2 ' h 0 0 0 0 0 0 7 e ;  
         r a m _ c e l l [           2 4 3 ]   =   3 2 ' h 0 0 0 0 0 0 0 0 ;  
         r a m _ c e l l [           2 4 4 ]   =   3 2 ' h 0 0 0 0 0 0 3 8 ;  
         r a m _ c e l l [           2 4 5 ]   =   3 2 ' h 0 0 0 0 0 0 1 6 ;  
         r a m _ c e l l [           2 4 6 ]   =   3 2 ' h 0 0 0 0 0 1 1 f ;  
         r a m _ c e l l [           2 4 7 ]   =   3 2 ' h 0 0 0 0 0 1 6 0 ;  
         r a m _ c e l l [           2 4 8 ]   =   3 2 ' h 0 0 0 0 0 1 a 1 ;  
         r a m _ c e l l [           2 4 9 ]   =   3 2 ' h 0 0 0 0 0 1 0 0 ;  
         r a m _ c e l l [           2 5 0 ]   =   3 2 ' h 0 0 0 0 0 0 b 5 ;  
         r a m _ c e l l [           2 5 1 ]   =   3 2 ' h 0 0 0 0 0 1 e b ;  
         r a m _ c e l l [           2 5 2 ]   =   3 2 ' h 0 0 0 0 0 0 5 8 ;  
         r a m _ c e l l [           2 5 3 ]   =   3 2 ' h 0 0 0 0 0 0 e 7 ;  
         r a m _ c e l l [           2 5 4 ]   =   3 2 ' h 0 0 0 0 0 1 9 f ;  
         r a m _ c e l l [           2 5 5 ]   =   3 2 ' h 0 0 0 0 0 0 4 9 ;  
         r a m _ c e l l [           2 5 6 ]   =   3 2 ' h 0 0 0 0 0 0 1 d ;  
         r a m _ c e l l [           2 5 7 ]   =   3 2 ' h 0 0 0 0 0 0 0 f ;  
         r a m _ c e l l [           2 5 8 ]   =   3 2 ' h 0 0 0 0 0 1 f 0 ;  
         r a m _ c e l l [           2 5 9 ]   =   3 2 ' h 0 0 0 0 0 0 3 e ;  
         r a m _ c e l l [           2 6 0 ]   =   3 2 ' h 0 0 0 0 0 0 e 8 ;  
         r a m _ c e l l [           2 6 1 ]   =   3 2 ' h 0 0 0 0 0 0 c f ;  
         r a m _ c e l l [           2 6 2 ]   =   3 2 ' h 0 0 0 0 0 1 4 4 ;  
         r a m _ c e l l [           2 6 3 ]   =   3 2 ' h 0 0 0 0 0 0 1 9 ;  
         r a m _ c e l l [           2 6 4 ]   =   3 2 ' h 0 0 0 0 0 1 2 5 ;  
         r a m _ c e l l [           2 6 5 ]   =   3 2 ' h 0 0 0 0 0 1 a 7 ;  
         r a m _ c e l l [           2 6 6 ]   =   3 2 ' h 0 0 0 0 0 1 2 d ;  
         r a m _ c e l l [           2 6 7 ]   =   3 2 ' h 0 0 0 0 0 1 3 f ;  
         r a m _ c e l l [           2 6 8 ]   =   3 2 ' h 0 0 0 0 0 1 3 d ;  
         r a m _ c e l l [           2 6 9 ]   =   3 2 ' h 0 0 0 0 0 0 a c ;  
         r a m _ c e l l [           2 7 0 ]   =   3 2 ' h 0 0 0 0 0 0 1 7 ;  
         r a m _ c e l l [           2 7 1 ]   =   3 2 ' h 0 0 0 0 0 1 c 8 ;  
         r a m _ c e l l [           2 7 2 ]   =   3 2 ' h 0 0 0 0 0 0 3 0 ;  
         r a m _ c e l l [           2 7 3 ]   =   3 2 ' h 0 0 0 0 0 0 4 f ;  
         r a m _ c e l l [           2 7 4 ]   =   3 2 ' h 0 0 0 0 0 1 5 0 ;  
         r a m _ c e l l [           2 7 5 ]   =   3 2 ' h 0 0 0 0 0 0 f 8 ;  
         r a m _ c e l l [           2 7 6 ]   =   3 2 ' h 0 0 0 0 0 1 c 6 ;  
         r a m _ c e l l [           2 7 7 ]   =   3 2 ' h 0 0 0 0 0 0 d 8 ;  
         r a m _ c e l l [           2 7 8 ]   =   3 2 ' h 0 0 0 0 0 0 2 a ;  
         r a m _ c e l l [           2 7 9 ]   =   3 2 ' h 0 0 0 0 0 1 3 e ;  
         r a m _ c e l l [           2 8 0 ]   =   3 2 ' h 0 0 0 0 0 0 8 f ;  
         r a m _ c e l l [           2 8 1 ]   =   3 2 ' h 0 0 0 0 0 0 f f ;  
         r a m _ c e l l [           2 8 2 ]   =   3 2 ' h 0 0 0 0 0 1 f b ;  
         r a m _ c e l l [           2 8 3 ]   =   3 2 ' h 0 0 0 0 0 0 2 1 ;  
         r a m _ c e l l [           2 8 4 ]   =   3 2 ' h 0 0 0 0 0 1 3 3 ;  
         r a m _ c e l l [           2 8 5 ]   =   3 2 ' h 0 0 0 0 0 1 4 b ;  
         r a m _ c e l l [           2 8 6 ]   =   3 2 ' h 0 0 0 0 0 1 a 4 ;  
         r a m _ c e l l [           2 8 7 ]   =   3 2 ' h 0 0 0 0 0 1 2 6 ;  
         r a m _ c e l l [           2 8 8 ]   =   3 2 ' h 0 0 0 0 0 1 3 b ;  
         r a m _ c e l l [           2 8 9 ]   =   3 2 ' h 0 0 0 0 0 1 5 a ;  
         r a m _ c e l l [           2 9 0 ]   =   3 2 ' h 0 0 0 0 0 1 b a ;  
         r a m _ c e l l [           2 9 1 ]   =   3 2 ' h 0 0 0 0 0 1 2 c ;  
         r a m _ c e l l [           2 9 2 ]   =   3 2 ' h 0 0 0 0 0 1 f 1 ;  
         r a m _ c e l l [           2 9 3 ]   =   3 2 ' h 0 0 0 0 0 0 b f ;  
         r a m _ c e l l [           2 9 4 ]   =   3 2 ' h 0 0 0 0 0 0 6 6 ;  
         r a m _ c e l l [           2 9 5 ]   =   3 2 ' h 0 0 0 0 0 0 8 b ;  
         r a m _ c e l l [           2 9 6 ]   =   3 2 ' h 0 0 0 0 0 0 f 2 ;  
         r a m _ c e l l [           2 9 7 ]   =   3 2 ' h 0 0 0 0 0 1 8 3 ;  
         r a m _ c e l l [           2 9 8 ]   =   3 2 ' h 0 0 0 0 0 1 c 5 ;  
         r a m _ c e l l [           2 9 9 ]   =   3 2 ' h 0 0 0 0 0 0 7 7 ;  
         r a m _ c e l l [           3 0 0 ]   =   3 2 ' h 0 0 0 0 0 1 a b ;  
         r a m _ c e l l [           3 0 1 ]   =   3 2 ' h 0 0 0 0 0 0 1 e ;  
         r a m _ c e l l [           3 0 2 ]   =   3 2 ' h 0 0 0 0 0 0 a 5 ;  
         r a m _ c e l l [           3 0 3 ]   =   3 2 ' h 0 0 0 0 0 1 9 0 ;  
         r a m _ c e l l [           3 0 4 ]   =   3 2 ' h 0 0 0 0 0 0 3 4 ;  
         r a m _ c e l l [           3 0 5 ]   =   3 2 ' h 0 0 0 0 0 1 7 3 ;  
         r a m _ c e l l [           3 0 6 ]   =   3 2 ' h 0 0 0 0 0 0 4 d ;  
         r a m _ c e l l [           3 0 7 ]   =   3 2 ' h 0 0 0 0 0 0 8 c ;  
         r a m _ c e l l [           3 0 8 ]   =   3 2 ' h 0 0 0 0 0 1 d 8 ;  
         r a m _ c e l l [           3 0 9 ]   =   3 2 ' h 0 0 0 0 0 0 5 2 ;  
         r a m _ c e l l [           3 1 0 ]   =   3 2 ' h 0 0 0 0 0 1 c 2 ;  
         r a m _ c e l l [           3 1 1 ]   =   3 2 ' h 0 0 0 0 0 1 8 b ;  
         r a m _ c e l l [           3 1 2 ]   =   3 2 ' h 0 0 0 0 0 0 9 8 ;  
         r a m _ c e l l [           3 1 3 ]   =   3 2 ' h 0 0 0 0 0 0 b 1 ;  
         r a m _ c e l l [           3 1 4 ]   =   3 2 ' h 0 0 0 0 0 1 6 7 ;  
         r a m _ c e l l [           3 1 5 ]   =   3 2 ' h 0 0 0 0 0 1 7 b ;  
         r a m _ c e l l [           3 1 6 ]   =   3 2 ' h 0 0 0 0 0 0 d 0 ;  
         r a m _ c e l l [           3 1 7 ]   =   3 2 ' h 0 0 0 0 0 0 5 3 ;  
         r a m _ c e l l [           3 1 8 ]   =   3 2 ' h 0 0 0 0 0 0 7 3 ;  
         r a m _ c e l l [           3 1 9 ]   =   3 2 ' h 0 0 0 0 0 0 f 3 ;  
         r a m _ c e l l [           3 2 0 ]   =   3 2 ' h 0 0 0 0 0 1 1 e ;  
         r a m _ c e l l [           3 2 1 ]   =   3 2 ' h 0 0 0 0 0 0 3 a ;  
         r a m _ c e l l [           3 2 2 ]   =   3 2 ' h 0 0 0 0 0 1 9 4 ;  
         r a m _ c e l l [           3 2 3 ]   =   3 2 ' h 0 0 0 0 0 1 3 1 ;  
         r a m _ c e l l [           3 2 4 ]   =   3 2 ' h 0 0 0 0 0 0 1 0 ;  
         r a m _ c e l l [           3 2 5 ]   =   3 2 ' h 0 0 0 0 0 0 b 2 ;  
         r a m _ c e l l [           3 2 6 ]   =   3 2 ' h 0 0 0 0 0 0 2 b ;  
         r a m _ c e l l [           3 2 7 ]   =   3 2 ' h 0 0 0 0 0 1 0 d ;  
         r a m _ c e l l [           3 2 8 ]   =   3 2 ' h 0 0 0 0 0 1 5 1 ;  
         r a m _ c e l l [           3 2 9 ]   =   3 2 ' h 0 0 0 0 0 1 8 4 ;  
         r a m _ c e l l [           3 3 0 ]   =   3 2 ' h 0 0 0 0 0 1 0 e ;  
         r a m _ c e l l [           3 3 1 ]   =   3 2 ' h 0 0 0 0 0 1 c 4 ;  
         r a m _ c e l l [           3 3 2 ]   =   3 2 ' h 0 0 0 0 0 1 c c ;  
         r a m _ c e l l [           3 3 3 ]   =   3 2 ' h 0 0 0 0 0 1 3 c ;  
         r a m _ c e l l [           3 3 4 ]   =   3 2 ' h 0 0 0 0 0 0 1 b ;  
         r a m _ c e l l [           3 3 5 ]   =   3 2 ' h 0 0 0 0 0 1 0 4 ;  
         r a m _ c e l l [           3 3 6 ]   =   3 2 ' h 0 0 0 0 0 0 7 4 ;  
         r a m _ c e l l [           3 3 7 ]   =   3 2 ' h 0 0 0 0 0 0 8 9 ;  
         r a m _ c e l l [           3 3 8 ]   =   3 2 ' h 0 0 0 0 0 1 5 b ;  
         r a m _ c e l l [           3 3 9 ]   =   3 2 ' h 0 0 0 0 0 1 9 6 ;  
         r a m _ c e l l [           3 4 0 ]   =   3 2 ' h 0 0 0 0 0 0 0 9 ;  
         r a m _ c e l l [           3 4 1 ]   =   3 2 ' h 0 0 0 0 0 0 c d ;  
         r a m _ c e l l [           3 4 2 ]   =   3 2 ' h 0 0 0 0 0 1 3 4 ;  
         r a m _ c e l l [           3 4 3 ]   =   3 2 ' h 0 0 0 0 0 0 a a ;  
         r a m _ c e l l [           3 4 4 ]   =   3 2 ' h 0 0 0 0 0 0 d c ;  
         r a m _ c e l l [           3 4 5 ]   =   3 2 ' h 0 0 0 0 0 1 c b ;  
         r a m _ c e l l [           3 4 6 ]   =   3 2 ' h 0 0 0 0 0 1 b 7 ;  
         r a m _ c e l l [           3 4 7 ]   =   3 2 ' h 0 0 0 0 0 0 5 b ;  
         r a m _ c e l l [           3 4 8 ]   =   3 2 ' h 0 0 0 0 0 1 7 2 ;  
         r a m _ c e l l [           3 4 9 ]   =   3 2 ' h 0 0 0 0 0 0 9 1 ;  
         r a m _ c e l l [           3 5 0 ]   =   3 2 ' h 0 0 0 0 0 1 1 6 ;  
         r a m _ c e l l [           3 5 1 ]   =   3 2 ' h 0 0 0 0 0 0 7 1 ;  
         r a m _ c e l l [           3 5 2 ]   =   3 2 ' h 0 0 0 0 0 1 6 8 ;  
         r a m _ c e l l [           3 5 3 ]   =   3 2 ' h 0 0 0 0 0 1 0 5 ;  
         r a m _ c e l l [           3 5 4 ]   =   3 2 ' h 0 0 0 0 0 0 3 6 ;  
         r a m _ c e l l [           3 5 5 ]   =   3 2 ' h 0 0 0 0 0 1 f a ;  
         r a m _ c e l l [           3 5 6 ]   =   3 2 ' h 0 0 0 0 0 1 7 4 ;  
         r a m _ c e l l [           3 5 7 ]   =   3 2 ' h 0 0 0 0 0 0 d d ;  
         r a m _ c e l l [           3 5 8 ]   =   3 2 ' h 0 0 0 0 0 1 d 7 ;  
         r a m _ c e l l [           3 5 9 ]   =   3 2 ' h 0 0 0 0 0 0 d 9 ;  
         r a m _ c e l l [           3 6 0 ]   =   3 2 ' h 0 0 0 0 0 0 c 9 ;  
         r a m _ c e l l [           3 6 1 ]   =   3 2 ' h 0 0 0 0 0 1 f f ;  
         r a m _ c e l l [           3 6 2 ]   =   3 2 ' h 0 0 0 0 0 0 5 d ;  
         r a m _ c e l l [           3 6 3 ]   =   3 2 ' h 0 0 0 0 0 1 8 d ;  
         r a m _ c e l l [           3 6 4 ]   =   3 2 ' h 0 0 0 0 0 1 7 1 ;  
         r a m _ c e l l [           3 6 5 ]   =   3 2 ' h 0 0 0 0 0 0 8 a ;  
         r a m _ c e l l [           3 6 6 ]   =   3 2 ' h 0 0 0 0 0 1 7 c ;  
         r a m _ c e l l [           3 6 7 ]   =   3 2 ' h 0 0 0 0 0 0 d 2 ;  
         r a m _ c e l l [           3 6 8 ]   =   3 2 ' h 0 0 0 0 0 0 c 4 ;  
         r a m _ c e l l [           3 6 9 ]   =   3 2 ' h 0 0 0 0 0 0 8 4 ;  
         r a m _ c e l l [           3 7 0 ]   =   3 2 ' h 0 0 0 0 0 0 2 2 ;  
         r a m _ c e l l [           3 7 1 ]   =   3 2 ' h 0 0 0 0 0 1 4 9 ;  
         r a m _ c e l l [           3 7 2 ]   =   3 2 ' h 0 0 0 0 0 0 5 a ;  
         r a m _ c e l l [           3 7 3 ]   =   3 2 ' h 0 0 0 0 0 0 9 4 ;  
         r a m _ c e l l [           3 7 4 ]   =   3 2 ' h 0 0 0 0 0 1 b c ;  
         r a m _ c e l l [           3 7 5 ]   =   3 2 ' h 0 0 0 0 0 0 c 3 ;  
         r a m _ c e l l [           3 7 6 ]   =   3 2 ' h 0 0 0 0 0 1 4 5 ;  
         r a m _ c e l l [           3 7 7 ]   =   3 2 ' h 0 0 0 0 0 0 c 1 ;  
         r a m _ c e l l [           3 7 8 ]   =   3 2 ' h 0 0 0 0 0 0 0 a ;  
         r a m _ c e l l [           3 7 9 ]   =   3 2 ' h 0 0 0 0 0 1 f e ;  
         r a m _ c e l l [           3 8 0 ]   =   3 2 ' h 0 0 0 0 0 0 b e ;  
         r a m _ c e l l [           3 8 1 ]   =   3 2 ' h 0 0 0 0 0 1 e c ;  
         r a m _ c e l l [           3 8 2 ]   =   3 2 ' h 0 0 0 0 0 0 f 4 ;  
         r a m _ c e l l [           3 8 3 ]   =   3 2 ' h 0 0 0 0 0 0 3 d ;  
         r a m _ c e l l [           3 8 4 ]   =   3 2 ' h 0 0 0 0 0 0 3 9 ;  
         r a m _ c e l l [           3 8 5 ]   =   3 2 ' h 0 0 0 0 0 0 8 8 ;  
         r a m _ c e l l [           3 8 6 ]   =   3 2 ' h 0 0 0 0 0 0 7 6 ;  
         r a m _ c e l l [           3 8 7 ]   =   3 2 ' h 0 0 0 0 0 0 4 5 ;  
         r a m _ c e l l [           3 8 8 ]   =   3 2 ' h 0 0 0 0 0 0 c 0 ;  
         r a m _ c e l l [           3 8 9 ]   =   3 2 ' h 0 0 0 0 0 0 f c ;  
         r a m _ c e l l [           3 9 0 ]   =   3 2 ' h 0 0 0 0 0 1 a 0 ;  
         r a m _ c e l l [           3 9 1 ]   =   3 2 ' h 0 0 0 0 0 1 9 2 ;  
         r a m _ c e l l [           3 9 2 ]   =   3 2 ' h 0 0 0 0 0 0 6 3 ;  
         r a m _ c e l l [           3 9 3 ]   =   3 2 ' h 0 0 0 0 0 1 d 5 ;  
         r a m _ c e l l [           3 9 4 ]   =   3 2 ' h 0 0 0 0 0 0 0 5 ;  
         r a m _ c e l l [           3 9 5 ]   =   3 2 ' h 0 0 0 0 0 1 a 3 ;  
         r a m _ c e l l [           3 9 6 ]   =   3 2 ' h 0 0 0 0 0 0 2 d ;  
         r a m _ c e l l [           3 9 7 ]   =   3 2 ' h 0 0 0 0 0 1 9 b ;  
         r a m _ c e l l [           3 9 8 ]   =   3 2 ' h 0 0 0 0 0 1 b 8 ;  
         r a m _ c e l l [           3 9 9 ]   =   3 2 ' h 0 0 0 0 0 0 c 6 ;  
         r a m _ c e l l [           4 0 0 ]   =   3 2 ' h 0 0 0 0 0 0 b c ;  
         r a m _ c e l l [           4 0 1 ]   =   3 2 ' h 0 0 0 0 0 1 b d ;  
         r a m _ c e l l [           4 0 2 ]   =   3 2 ' h 0 0 0 0 0 1 7 e ;  
         r a m _ c e l l [           4 0 3 ]   =   3 2 ' h 0 0 0 0 0 1 4 a ;  
         r a m _ c e l l [           4 0 4 ]   =   3 2 ' h 0 0 0 0 0 0 6 9 ;  
         r a m _ c e l l [           4 0 5 ]   =   3 2 ' h 0 0 0 0 0 1 b 1 ;  
         r a m _ c e l l [           4 0 6 ]   =   3 2 ' h 0 0 0 0 0 1 0 1 ;  
         r a m _ c e l l [           4 0 7 ]   =   3 2 ' h 0 0 0 0 0 1 0 f ;  
         r a m _ c e l l [           4 0 8 ]   =   3 2 ' h 0 0 0 0 0 0 5 7 ;  
         r a m _ c e l l [           4 0 9 ]   =   3 2 ' h 0 0 0 0 0 1 b 5 ;  
         r a m _ c e l l [           4 1 0 ]   =   3 2 ' h 0 0 0 0 0 1 2 7 ;  
         r a m _ c e l l [           4 1 1 ]   =   3 2 ' h 0 0 0 0 0 1 8 7 ;  
         r a m _ c e l l [           4 1 2 ]   =   3 2 ' h 0 0 0 0 0 0 8 6 ;  
         r a m _ c e l l [           4 1 3 ]   =   3 2 ' h 0 0 0 0 0 0 6 e ;  
         r a m _ c e l l [           4 1 4 ]   =   3 2 ' h 0 0 0 0 0 0 7 d ;  
         r a m _ c e l l [           4 1 5 ]   =   3 2 ' h 0 0 0 0 0 1 9 8 ;  
         r a m _ c e l l [           4 1 6 ]   =   3 2 ' h 0 0 0 0 0 1 b 6 ;  
         r a m _ c e l l [           4 1 7 ]   =   3 2 ' h 0 0 0 0 0 0 2 4 ;  
         r a m _ c e l l [           4 1 8 ]   =   3 2 ' h 0 0 0 0 0 0 9 a ;  
         r a m _ c e l l [           4 1 9 ]   =   3 2 ' h 0 0 0 0 0 1 a 9 ;  
         r a m _ c e l l [           4 2 0 ]   =   3 2 ' h 0 0 0 0 0 0 6 4 ;  
         r a m _ c e l l [           4 2 1 ]   =   3 2 ' h 0 0 0 0 0 0 3 f ;  
         r a m _ c e l l [           4 2 2 ]   =   3 2 ' h 0 0 0 0 0 1 1 b ;  
         r a m _ c e l l [           4 2 3 ]   =   3 2 ' h 0 0 0 0 0 1 a 2 ;  
         r a m _ c e l l [           4 2 4 ]   =   3 2 ' h 0 0 0 0 0 1 9 c ;  
         r a m _ c e l l [           4 2 5 ]   =   3 2 ' h 0 0 0 0 0 1 5 7 ;  
         r a m _ c e l l [           4 2 6 ]   =   3 2 ' h 0 0 0 0 0 0 4 3 ;  
         r a m _ c e l l [           4 2 7 ]   =   3 2 ' h 0 0 0 0 0 0 e f ;  
         r a m _ c e l l [           4 2 8 ]   =   3 2 ' h 0 0 0 0 0 0 4 0 ;  
         r a m _ c e l l [           4 2 9 ]   =   3 2 ' h 0 0 0 0 0 0 3 b ;  
         r a m _ c e l l [           4 3 0 ]   =   3 2 ' h 0 0 0 0 0 0 f 0 ;  
         r a m _ c e l l [           4 3 1 ]   =   3 2 ' h 0 0 0 0 0 1 d 6 ;  
         r a m _ c e l l [           4 3 2 ]   =   3 2 ' h 0 0 0 0 0 1 6 c ;  
         r a m _ c e l l [           4 3 3 ]   =   3 2 ' h 0 0 0 0 0 0 2 8 ;  
         r a m _ c e l l [           4 3 4 ]   =   3 2 ' h 0 0 0 0 0 0 a 7 ;  
         r a m _ c e l l [           4 3 5 ]   =   3 2 ' h 0 0 0 0 0 1 6 9 ;  
         r a m _ c e l l [           4 3 6 ]   =   3 2 ' h 0 0 0 0 0 1 d d ;  
         r a m _ c e l l [           4 3 7 ]   =   3 2 ' h 0 0 0 0 0 0 7 f ;  
         r a m _ c e l l [           4 3 8 ]   =   3 2 ' h 0 0 0 0 0 0 d 3 ;  
         r a m _ c e l l [           4 3 9 ]   =   3 2 ' h 0 0 0 0 0 1 2 b ;  
         r a m _ c e l l [           4 4 0 ]   =   3 2 ' h 0 0 0 0 0 0 1 a ;  
         r a m _ c e l l [           4 4 1 ]   =   3 2 ' h 0 0 0 0 0 0 c b ;  
         r a m _ c e l l [           4 4 2 ]   =   3 2 ' h 0 0 0 0 0 0 4 6 ;  
         r a m _ c e l l [           4 4 3 ]   =   3 2 ' h 0 0 0 0 0 0 a 2 ;  
         r a m _ c e l l [           4 4 4 ]   =   3 2 ' h 0 0 0 0 0 1 d c ;  
         r a m _ c e l l [           4 4 5 ]   =   3 2 ' h 0 0 0 0 0 0 9 d ;  
         r a m _ c e l l [           4 4 6 ]   =   3 2 ' h 0 0 0 0 0 0 f e ;  
         r a m _ c e l l [           4 4 7 ]   =   3 2 ' h 0 0 0 0 0 0 a 1 ;  
         r a m _ c e l l [           4 4 8 ]   =   3 2 ' h 0 0 0 0 0 1 d 3 ;  
         r a m _ c e l l [           4 4 9 ]   =   3 2 ' h 0 0 0 0 0 0 a 3 ;  
         r a m _ c e l l [           4 5 0 ]   =   3 2 ' h 0 0 0 0 0 1 6 1 ;  
         r a m _ c e l l [           4 5 1 ]   =   3 2 ' h 0 0 0 0 0 0 d e ;  
         r a m _ c e l l [           4 5 2 ]   =   3 2 ' h 0 0 0 0 0 1 8 8 ;  
         r a m _ c e l l [           4 5 3 ]   =   3 2 ' h 0 0 0 0 0 1 f 7 ;  
         r a m _ c e l l [           4 5 4 ]   =   3 2 ' h 0 0 0 0 0 1 5 2 ;  
         r a m _ c e l l [           4 5 5 ]   =   3 2 ' h 0 0 0 0 0 1 3 9 ;  
         r a m _ c e l l [           4 5 6 ]   =   3 2 ' h 0 0 0 0 0 0 7 c ;  
         r a m _ c e l l [           4 5 7 ]   =   3 2 ' h 0 0 0 0 0 0 2 3 ;  
         r a m _ c e l l [           4 5 8 ]   =   3 2 ' h 0 0 0 0 0 1 3 a ;  
         r a m _ c e l l [           4 5 9 ]   =   3 2 ' h 0 0 0 0 0 1 c f ;  
         r a m _ c e l l [           4 6 0 ]   =   3 2 ' h 0 0 0 0 0 1 e e ;  
         r a m _ c e l l [           4 6 1 ]   =   3 2 ' h 0 0 0 0 0 1 4 6 ;  
         r a m _ c e l l [           4 6 2 ]   =   3 2 ' h 0 0 0 0 0 0 d 6 ;  
         r a m _ c e l l [           4 6 3 ]   =   3 2 ' h 0 0 0 0 0 1 5 3 ;  
         r a m _ c e l l [           4 6 4 ]   =   3 2 ' h 0 0 0 0 0 0 d a ;  
         r a m _ c e l l [           4 6 5 ]   =   3 2 ' h 0 0 0 0 0 1 d 4 ;  
         r a m _ c e l l [           4 6 6 ]   =   3 2 ' h 0 0 0 0 0 0 7 b ;  
         r a m _ c e l l [           4 6 7 ]   =   3 2 ' h 0 0 0 0 0 0 8 0 ;  
         r a m _ c e l l [           4 6 8 ]   =   3 2 ' h 0 0 0 0 0 0 e 2 ;  
         r a m _ c e l l [           4 6 9 ]   =   3 2 ' h 0 0 0 0 0 0 e 4 ;  
         r a m _ c e l l [           4 7 0 ]   =   3 2 ' h 0 0 0 0 0 0 0 7 ;  
         r a m _ c e l l [           4 7 1 ]   =   3 2 ' h 0 0 0 0 0 0 9 5 ;  
         r a m _ c e l l [           4 7 2 ]   =   3 2 ' h 0 0 0 0 0 1 6 e ;  
         r a m _ c e l l [           4 7 3 ]   =   3 2 ' h 0 0 0 0 0 0 b 4 ;  
         r a m _ c e l l [           4 7 4 ]   =   3 2 ' h 0 0 0 0 0 0 9 0 ;  
         r a m _ c e l l [           4 7 5 ]   =   3 2 ' h 0 0 0 0 0 1 4 c ;  
         r a m _ c e l l [           4 7 6 ]   =   3 2 ' h 0 0 0 0 0 0 0 2 ;  
         r a m _ c e l l [           4 7 7 ]   =   3 2 ' h 0 0 0 0 0 0 e 0 ;  
         r a m _ c e l l [           4 7 8 ]   =   3 2 ' h 0 0 0 0 0 0 c 8 ;  
         r a m _ c e l l [           4 7 9 ]   =   3 2 ' h 0 0 0 0 0 1 1 c ;  
         r a m _ c e l l [           4 8 0 ]   =   3 2 ' h 0 0 0 0 0 0 0 8 ;  
         r a m _ c e l l [           4 8 1 ]   =   3 2 ' h 0 0 0 0 0 0 6 a ;  
         r a m _ c e l l [           4 8 2 ]   =   3 2 ' h 0 0 0 0 0 1 7 6 ;  
         r a m _ c e l l [           4 8 3 ]   =   3 2 ' h 0 0 0 0 0 1 1 d ;  
         r a m _ c e l l [           4 8 4 ]   =   3 2 ' h 0 0 0 0 0 1 e 4 ;  
         r a m _ c e l l [           4 8 5 ]   =   3 2 ' h 0 0 0 0 0 1 d a ;  
         r a m _ c e l l [           4 8 6 ]   =   3 2 ' h 0 0 0 0 0 1 7 a ;  
         r a m _ c e l l [           4 8 7 ]   =   3 2 ' h 0 0 0 0 0 1 e 1 ;  
         r a m _ c e l l [           4 8 8 ]   =   3 2 ' h 0 0 0 0 0 0 6 d ;  
         r a m _ c e l l [           4 8 9 ]   =   3 2 ' h 0 0 0 0 0 0 1 3 ;  
         r a m _ c e l l [           4 9 0 ]   =   3 2 ' h 0 0 0 0 0 0 e 9 ;  
         r a m _ c e l l [           4 9 1 ]   =   3 2 ' h 0 0 0 0 0 1 1 7 ;  
         r a m _ c e l l [           4 9 2 ]   =   3 2 ' h 0 0 0 0 0 1 f 4 ;  
         r a m _ c e l l [           4 9 3 ]   =   3 2 ' h 0 0 0 0 0 1 7 7 ;  
         r a m _ c e l l [           4 9 4 ]   =   3 2 ' h 0 0 0 0 0 0 5 f ;  
         r a m _ c e l l [           4 9 5 ]   =   3 2 ' h 0 0 0 0 0 1 3 0 ;  
         r a m _ c e l l [           4 9 6 ]   =   3 2 ' h 0 0 0 0 0 0 a 0 ;  
         r a m _ c e l l [           4 9 7 ]   =   3 2 ' h 0 0 0 0 0 0 e 1 ;  
         r a m _ c e l l [           4 9 8 ]   =   3 2 ' h 0 0 0 0 0 1 2 9 ;  
         r a m _ c e l l [           4 9 9 ]   =   3 2 ' h 0 0 0 0 0 0 f 1 ;  
         r a m _ c e l l [           5 0 0 ]   =   3 2 ' h 0 0 0 0 0 1 7 d ;  
         r a m _ c e l l [           5 0 1 ]   =   3 2 ' h 0 0 0 0 0 1 0 c ;  
         r a m _ c e l l [           5 0 2 ]   =   3 2 ' h 0 0 0 0 0 1 f d ;  
         r a m _ c e l l [           5 0 3 ]   =   3 2 ' h 0 0 0 0 0 0 a d ;  
         r a m _ c e l l [           5 0 4 ]   =   3 2 ' h 0 0 0 0 0 0 8 e ;  
         r a m _ c e l l [           5 0 5 ]   =   3 2 ' h 0 0 0 0 0 1 c e ;  
         r a m _ c e l l [           5 0 6 ]   =   3 2 ' h 0 0 0 0 0 1 2 3 ;  
         r a m _ c e l l [           5 0 7 ]   =   3 2 ' h 0 0 0 0 0 0 9 9 ;  
         r a m _ c e l l [           5 0 8 ]   =   3 2 ' h 0 0 0 0 0 1 b e ;  
         r a m _ c e l l [           5 0 9 ]   =   3 2 ' h 0 0 0 0 0 0 9 6 ;  
         r a m _ c e l l [           5 1 0 ]   =   3 2 ' h 0 0 0 0 0 0 4 1 ;  
         r a m _ c e l l [           5 1 1 ]   =   3 2 ' h 0 0 0 0 0 1 8 1 ;  
 e n d  
  
 e n d m o d u l e  
  
 