
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    ram_cell[       0] = 32'h000001ac;
    ram_cell[       1] = 32'h000000d0;
    ram_cell[       2] = 32'h00000067;
    ram_cell[       3] = 32'h000000ff;
    ram_cell[       4] = 32'h0000012f;
    ram_cell[       5] = 32'h000001b6;
    ram_cell[       6] = 32'h000000ed;
    ram_cell[       7] = 32'h000001ef;
    ram_cell[       8] = 32'h00000102;
    ram_cell[       9] = 32'h00000045;
    ram_cell[      10] = 32'h00000028;
    ram_cell[      11] = 32'h0000000c;
    ram_cell[      12] = 32'h00000078;
    ram_cell[      13] = 32'h00000072;
    ram_cell[      14] = 32'h000001b0;
    ram_cell[      15] = 32'h000001ad;
    ram_cell[      16] = 32'h000000e8;
    ram_cell[      17] = 32'h00000154;
    ram_cell[      18] = 32'h000000cc;
    ram_cell[      19] = 32'h000000df;
    ram_cell[      20] = 32'h0000004e;
    ram_cell[      21] = 32'h000000be;
    ram_cell[      22] = 32'h000000cb;
    ram_cell[      23] = 32'h00000074;
    ram_cell[      24] = 32'h000000fb;
    ram_cell[      25] = 32'h000000db;
    ram_cell[      26] = 32'h00000033;
    ram_cell[      27] = 32'h0000012a;
    ram_cell[      28] = 32'h000000cf;
    ram_cell[      29] = 32'h000000f1;
    ram_cell[      30] = 32'h00000129;
    ram_cell[      31] = 32'h0000016f;
    ram_cell[      32] = 32'h000000b5;
    ram_cell[      33] = 32'h00000092;
    ram_cell[      34] = 32'h000001a3;
    ram_cell[      35] = 32'h000001b2;
    ram_cell[      36] = 32'h00000047;
    ram_cell[      37] = 32'h00000147;
    ram_cell[      38] = 32'h00000149;
    ram_cell[      39] = 32'h00000188;
    ram_cell[      40] = 32'h00000039;
    ram_cell[      41] = 32'h000000e0;
    ram_cell[      42] = 32'h00000187;
    ram_cell[      43] = 32'h00000166;
    ram_cell[      44] = 32'h000001bc;
    ram_cell[      45] = 32'h000000e7;
    ram_cell[      46] = 32'h000000f7;
    ram_cell[      47] = 32'h00000029;
    ram_cell[      48] = 32'h0000019d;
    ram_cell[      49] = 32'h0000005c;
    ram_cell[      50] = 32'h000001c1;
    ram_cell[      51] = 32'h000000ef;
    ram_cell[      52] = 32'h0000000f;
    ram_cell[      53] = 32'h000000f8;
    ram_cell[      54] = 32'h000000b8;
    ram_cell[      55] = 32'h00000038;
    ram_cell[      56] = 32'h00000097;
    ram_cell[      57] = 32'h00000043;
    ram_cell[      58] = 32'h000000ec;
    ram_cell[      59] = 32'h00000109;
    ram_cell[      60] = 32'h00000006;
    ram_cell[      61] = 32'h000001c6;
    ram_cell[      62] = 32'h000001bd;
    ram_cell[      63] = 32'h00000118;
    ram_cell[      64] = 32'h000001a9;
    ram_cell[      65] = 32'h0000003a;
    ram_cell[      66] = 32'h00000019;
    ram_cell[      67] = 32'h00000059;
    ram_cell[      68] = 32'h000001e0;
    ram_cell[      69] = 32'h000001d4;
    ram_cell[      70] = 32'h000000c9;
    ram_cell[      71] = 32'h000000d6;
    ram_cell[      72] = 32'h000000d2;
    ram_cell[      73] = 32'h00000191;
    ram_cell[      74] = 32'h0000013f;
    ram_cell[      75] = 32'h0000008e;
    ram_cell[      76] = 32'h000001ee;
    ram_cell[      77] = 32'h00000060;
    ram_cell[      78] = 32'h00000108;
    ram_cell[      79] = 32'h000000d3;
    ram_cell[      80] = 32'h0000006e;
    ram_cell[      81] = 32'h000000a0;
    ram_cell[      82] = 32'h000001f0;
    ram_cell[      83] = 32'h00000178;
    ram_cell[      84] = 32'h00000023;
    ram_cell[      85] = 32'h000000f3;
    ram_cell[      86] = 32'h000001a1;
    ram_cell[      87] = 32'h00000015;
    ram_cell[      88] = 32'h0000007b;
    ram_cell[      89] = 32'h000001b5;
    ram_cell[      90] = 32'h00000195;
    ram_cell[      91] = 32'h00000073;
    ram_cell[      92] = 32'h0000001b;
    ram_cell[      93] = 32'h0000007e;
    ram_cell[      94] = 32'h000001db;
    ram_cell[      95] = 32'h0000009c;
    ram_cell[      96] = 32'h0000007a;
    ram_cell[      97] = 32'h000000ca;
    ram_cell[      98] = 32'h000001eb;
    ram_cell[      99] = 32'h0000008f;
    ram_cell[     100] = 32'h0000009f;
    ram_cell[     101] = 32'h0000001d;
    ram_cell[     102] = 32'h0000019e;
    ram_cell[     103] = 32'h000000f2;
    ram_cell[     104] = 32'h00000116;
    ram_cell[     105] = 32'h000000da;
    ram_cell[     106] = 32'h000001c8;
    ram_cell[     107] = 32'h000001bf;
    ram_cell[     108] = 32'h00000130;
    ram_cell[     109] = 32'h000001ab;
    ram_cell[     110] = 32'h0000012d;
    ram_cell[     111] = 32'h00000125;
    ram_cell[     112] = 32'h00000064;
    ram_cell[     113] = 32'h0000001a;
    ram_cell[     114] = 32'h00000182;
    ram_cell[     115] = 32'h000000f4;
    ram_cell[     116] = 32'h00000139;
    ram_cell[     117] = 32'h000000fd;
    ram_cell[     118] = 32'h0000018e;
    ram_cell[     119] = 32'h0000015d;
    ram_cell[     120] = 32'h00000070;
    ram_cell[     121] = 32'h000000c7;
    ram_cell[     122] = 32'h0000002b;
    ram_cell[     123] = 32'h000001c2;
    ram_cell[     124] = 32'h00000145;
    ram_cell[     125] = 32'h0000007c;
    ram_cell[     126] = 32'h000001fd;
    ram_cell[     127] = 32'h000001e8;
    ram_cell[     128] = 32'h0000009a;
    ram_cell[     129] = 32'h00000197;
    ram_cell[     130] = 32'h00000194;
    ram_cell[     131] = 32'h00000111;
    ram_cell[     132] = 32'h00000050;
    ram_cell[     133] = 32'h00000176;
    ram_cell[     134] = 32'h000000aa;
    ram_cell[     135] = 32'h000001b4;
    ram_cell[     136] = 32'h000000e4;
    ram_cell[     137] = 32'h0000014b;
    ram_cell[     138] = 32'h000001f4;
    ram_cell[     139] = 32'h000000ce;
    ram_cell[     140] = 32'h00000146;
    ram_cell[     141] = 32'h00000104;
    ram_cell[     142] = 32'h00000017;
    ram_cell[     143] = 32'h00000168;
    ram_cell[     144] = 32'h00000003;
    ram_cell[     145] = 32'h00000012;
    ram_cell[     146] = 32'h00000071;
    ram_cell[     147] = 32'h00000052;
    ram_cell[     148] = 32'h0000009e;
    ram_cell[     149] = 32'h000000b6;
    ram_cell[     150] = 32'h00000141;
    ram_cell[     151] = 32'h00000009;
    ram_cell[     152] = 32'h00000170;
    ram_cell[     153] = 32'h000001f2;
    ram_cell[     154] = 32'h00000077;
    ram_cell[     155] = 32'h000000f9;
    ram_cell[     156] = 32'h00000075;
    ram_cell[     157] = 32'h00000153;
    ram_cell[     158] = 32'h00000044;
    ram_cell[     159] = 32'h000000a2;
    ram_cell[     160] = 32'h0000005e;
    ram_cell[     161] = 32'h000001cf;
    ram_cell[     162] = 32'h000001da;
    ram_cell[     163] = 32'h0000019c;
    ram_cell[     164] = 32'h00000048;
    ram_cell[     165] = 32'h00000113;
    ram_cell[     166] = 32'h00000081;
    ram_cell[     167] = 32'h0000000d;
    ram_cell[     168] = 32'h0000015a;
    ram_cell[     169] = 32'h00000098;
    ram_cell[     170] = 32'h00000087;
    ram_cell[     171] = 32'h00000193;
    ram_cell[     172] = 32'h00000156;
    ram_cell[     173] = 32'h00000080;
    ram_cell[     174] = 32'h000000f5;
    ram_cell[     175] = 32'h000000a7;
    ram_cell[     176] = 32'h000001de;
    ram_cell[     177] = 32'h0000012b;
    ram_cell[     178] = 32'h000000fc;
    ram_cell[     179] = 32'h0000017b;
    ram_cell[     180] = 32'h00000105;
    ram_cell[     181] = 32'h0000012e;
    ram_cell[     182] = 32'h000000b7;
    ram_cell[     183] = 32'h00000107;
    ram_cell[     184] = 32'h000000b3;
    ram_cell[     185] = 32'h0000001f;
    ram_cell[     186] = 32'h0000004d;
    ram_cell[     187] = 32'h00000094;
    ram_cell[     188] = 32'h00000083;
    ram_cell[     189] = 32'h00000167;
    ram_cell[     190] = 32'h000001a7;
    ram_cell[     191] = 32'h0000010a;
    ram_cell[     192] = 32'h000000e6;
    ram_cell[     193] = 32'h000000b1;
    ram_cell[     194] = 32'h000000dc;
    ram_cell[     195] = 32'h000001e6;
    ram_cell[     196] = 32'h00000138;
    ram_cell[     197] = 32'h00000171;
    ram_cell[     198] = 32'h000001df;
    ram_cell[     199] = 32'h00000016;
    ram_cell[     200] = 32'h000000b0;
    ram_cell[     201] = 32'h00000008;
    ram_cell[     202] = 32'h0000018f;
    ram_cell[     203] = 32'h0000006b;
    ram_cell[     204] = 32'h000000a6;
    ram_cell[     205] = 32'h0000016a;
    ram_cell[     206] = 32'h00000123;
    ram_cell[     207] = 32'h00000054;
    ram_cell[     208] = 32'h0000006c;
    ram_cell[     209] = 32'h0000014c;
    ram_cell[     210] = 32'h000000bc;
    ram_cell[     211] = 32'h0000000a;
    ram_cell[     212] = 32'h000001e3;
    ram_cell[     213] = 32'h00000175;
    ram_cell[     214] = 32'h00000106;
    ram_cell[     215] = 32'h000000b2;
    ram_cell[     216] = 32'h0000004f;
    ram_cell[     217] = 32'h000000c6;
    ram_cell[     218] = 32'h000001f8;
    ram_cell[     219] = 32'h00000110;
    ram_cell[     220] = 32'h00000088;
    ram_cell[     221] = 32'h00000036;
    ram_cell[     222] = 32'h00000062;
    ram_cell[     223] = 32'h000001d9;
    ram_cell[     224] = 32'h00000152;
    ram_cell[     225] = 32'h000000ae;
    ram_cell[     226] = 32'h000000eb;
    ram_cell[     227] = 32'h00000190;
    ram_cell[     228] = 32'h0000010e;
    ram_cell[     229] = 32'h000000d9;
    ram_cell[     230] = 32'h0000009b;
    ram_cell[     231] = 32'h0000008c;
    ram_cell[     232] = 32'h0000015f;
    ram_cell[     233] = 32'h000000f0;
    ram_cell[     234] = 32'h000000d8;
    ram_cell[     235] = 32'h00000189;
    ram_cell[     236] = 32'h00000132;
    ram_cell[     237] = 32'h0000005f;
    ram_cell[     238] = 32'h000001c3;
    ram_cell[     239] = 32'h000000d4;
    ram_cell[     240] = 32'h000000f6;
    ram_cell[     241] = 32'h000001cd;
    ram_cell[     242] = 32'h000000d1;
    ram_cell[     243] = 32'h00000049;
    ram_cell[     244] = 32'h0000015e;
    ram_cell[     245] = 32'h00000165;
    ram_cell[     246] = 32'h00000024;
    ram_cell[     247] = 32'h0000010d;
    ram_cell[     248] = 32'h00000022;
    ram_cell[     249] = 32'h0000015b;
    ram_cell[     250] = 32'h0000003c;
    ram_cell[     251] = 32'h00000084;
    ram_cell[     252] = 32'h000001dd;
    ram_cell[     253] = 32'h00000005;
    ram_cell[     254] = 32'h00000096;
    ram_cell[     255] = 32'h00000007;
    ram_cell[     256] = 32'h0000010b;
    ram_cell[     257] = 32'h000001d7;
    ram_cell[     258] = 32'h000001f6;
    ram_cell[     259] = 32'h00000164;
    ram_cell[     260] = 32'h00000093;
    ram_cell[     261] = 32'h0000003b;
    ram_cell[     262] = 32'h000000a3;
    ram_cell[     263] = 32'h0000010c;
    ram_cell[     264] = 32'h0000018a;
    ram_cell[     265] = 32'h00000095;
    ram_cell[     266] = 32'h00000056;
    ram_cell[     267] = 32'h00000032;
    ram_cell[     268] = 32'h000000af;
    ram_cell[     269] = 32'h000001b8;
    ram_cell[     270] = 32'h00000160;
    ram_cell[     271] = 32'h000000e1;
    ram_cell[     272] = 32'h00000199;
    ram_cell[     273] = 32'h00000076;
    ram_cell[     274] = 32'h0000008d;
    ram_cell[     275] = 32'h00000173;
    ram_cell[     276] = 32'h000001ae;
    ram_cell[     277] = 32'h0000003e;
    ram_cell[     278] = 32'h000000ba;
    ram_cell[     279] = 32'h0000011e;
    ram_cell[     280] = 32'h0000017f;
    ram_cell[     281] = 32'h000001ff;
    ram_cell[     282] = 32'h0000015c;
    ram_cell[     283] = 32'h000001a0;
    ram_cell[     284] = 32'h0000018c;
    ram_cell[     285] = 32'h00000014;
    ram_cell[     286] = 32'h000000c8;
    ram_cell[     287] = 32'h00000158;
    ram_cell[     288] = 32'h000001d0;
    ram_cell[     289] = 32'h00000172;
    ram_cell[     290] = 32'h0000010f;
    ram_cell[     291] = 32'h00000061;
    ram_cell[     292] = 32'h000000d7;
    ram_cell[     293] = 32'h000001f7;
    ram_cell[     294] = 32'h000001a4;
    ram_cell[     295] = 32'h0000013d;
    ram_cell[     296] = 32'h00000085;
    ram_cell[     297] = 32'h00000068;
    ram_cell[     298] = 32'h0000014f;
    ram_cell[     299] = 32'h00000128;
    ram_cell[     300] = 32'h00000037;
    ram_cell[     301] = 32'h000001ca;
    ram_cell[     302] = 32'h00000163;
    ram_cell[     303] = 32'h00000196;
    ram_cell[     304] = 32'h000001f1;
    ram_cell[     305] = 32'h0000005d;
    ram_cell[     306] = 32'h0000011f;
    ram_cell[     307] = 32'h000001c7;
    ram_cell[     308] = 32'h0000016e;
    ram_cell[     309] = 32'h00000140;
    ram_cell[     310] = 32'h00000020;
    ram_cell[     311] = 32'h00000063;
    ram_cell[     312] = 32'h00000121;
    ram_cell[     313] = 32'h00000134;
    ram_cell[     314] = 32'h00000013;
    ram_cell[     315] = 32'h0000003d;
    ram_cell[     316] = 32'h0000004c;
    ram_cell[     317] = 32'h00000089;
    ram_cell[     318] = 32'h00000030;
    ram_cell[     319] = 32'h000000c3;
    ram_cell[     320] = 32'h000001b1;
    ram_cell[     321] = 32'h0000018d;
    ram_cell[     322] = 32'h0000019a;
    ram_cell[     323] = 32'h000001cb;
    ram_cell[     324] = 32'h00000112;
    ram_cell[     325] = 32'h000000c4;
    ram_cell[     326] = 32'h00000192;
    ram_cell[     327] = 32'h000001c0;
    ram_cell[     328] = 32'h000001e2;
    ram_cell[     329] = 32'h000001fb;
    ram_cell[     330] = 32'h00000091;
    ram_cell[     331] = 32'h00000058;
    ram_cell[     332] = 32'h00000155;
    ram_cell[     333] = 32'h00000103;
    ram_cell[     334] = 32'h0000019b;
    ram_cell[     335] = 32'h0000000e;
    ram_cell[     336] = 32'h00000181;
    ram_cell[     337] = 32'h000001d3;
    ram_cell[     338] = 32'h0000008a;
    ram_cell[     339] = 32'h00000148;
    ram_cell[     340] = 32'h000001ec;
    ram_cell[     341] = 32'h0000011b;
    ram_cell[     342] = 32'h00000114;
    ram_cell[     343] = 32'h0000008b;
    ram_cell[     344] = 32'h000000c5;
    ram_cell[     345] = 32'h000000ab;
    ram_cell[     346] = 32'h0000002d;
    ram_cell[     347] = 32'h0000019f;
    ram_cell[     348] = 32'h000000a8;
    ram_cell[     349] = 32'h00000151;
    ram_cell[     350] = 32'h000000fa;
    ram_cell[     351] = 32'h000001d8;
    ram_cell[     352] = 32'h00000180;
    ram_cell[     353] = 32'h00000198;
    ram_cell[     354] = 32'h00000010;
    ram_cell[     355] = 32'h000001e1;
    ram_cell[     356] = 32'h000001d6;
    ram_cell[     357] = 32'h000000e3;
    ram_cell[     358] = 32'h00000053;
    ram_cell[     359] = 32'h0000005a;
    ram_cell[     360] = 32'h000001d1;
    ram_cell[     361] = 32'h00000131;
    ram_cell[     362] = 32'h000001c5;
    ram_cell[     363] = 32'h00000000;
    ram_cell[     364] = 32'h000000fe;
    ram_cell[     365] = 32'h000001a2;
    ram_cell[     366] = 32'h0000006a;
    ram_cell[     367] = 32'h000001e9;
    ram_cell[     368] = 32'h0000002a;
    ram_cell[     369] = 32'h00000144;
    ram_cell[     370] = 32'h000000c0;
    ram_cell[     371] = 32'h0000006f;
    ram_cell[     372] = 32'h0000016d;
    ram_cell[     373] = 32'h000000cd;
    ram_cell[     374] = 32'h00000143;
    ram_cell[     375] = 32'h000000e9;
    ram_cell[     376] = 32'h000000a4;
    ram_cell[     377] = 32'h000001fe;
    ram_cell[     378] = 32'h0000017c;
    ram_cell[     379] = 32'h00000120;
    ram_cell[     380] = 32'h000000b9;
    ram_cell[     381] = 32'h00000115;
    ram_cell[     382] = 32'h000000dd;
    ram_cell[     383] = 32'h000001b3;
    ram_cell[     384] = 32'h00000122;
    ram_cell[     385] = 32'h000001e4;
    ram_cell[     386] = 32'h000000de;
    ram_cell[     387] = 32'h00000161;
    ram_cell[     388] = 32'h000001ea;
    ram_cell[     389] = 32'h000000bb;
    ram_cell[     390] = 32'h000001f9;
    ram_cell[     391] = 32'h0000013e;
    ram_cell[     392] = 32'h000001a8;
    ram_cell[     393] = 32'h00000179;
    ram_cell[     394] = 32'h00000169;
    ram_cell[     395] = 32'h000001fa;
    ram_cell[     396] = 32'h00000066;
    ram_cell[     397] = 32'h00000034;
    ram_cell[     398] = 32'h000000ac;
    ram_cell[     399] = 32'h00000031;
    ram_cell[     400] = 32'h00000117;
    ram_cell[     401] = 32'h000001b9;
    ram_cell[     402] = 32'h000001a5;
    ram_cell[     403] = 32'h000001dc;
    ram_cell[     404] = 32'h00000042;
    ram_cell[     405] = 32'h000001e7;
    ram_cell[     406] = 32'h00000026;
    ram_cell[     407] = 32'h0000009d;
    ram_cell[     408] = 32'h0000014a;
    ram_cell[     409] = 32'h0000001c;
    ram_cell[     410] = 32'h00000011;
    ram_cell[     411] = 32'h00000018;
    ram_cell[     412] = 32'h00000101;
    ram_cell[     413] = 32'h00000055;
    ram_cell[     414] = 32'h000001b7;
    ram_cell[     415] = 32'h00000186;
    ram_cell[     416] = 32'h00000133;
    ram_cell[     417] = 32'h00000021;
    ram_cell[     418] = 32'h0000016b;
    ram_cell[     419] = 32'h0000011a;
    ram_cell[     420] = 32'h0000007f;
    ram_cell[     421] = 32'h00000027;
    ram_cell[     422] = 32'h0000003f;
    ram_cell[     423] = 32'h0000013a;
    ram_cell[     424] = 32'h0000017d;
    ram_cell[     425] = 32'h00000035;
    ram_cell[     426] = 32'h0000005b;
    ram_cell[     427] = 32'h0000007d;
    ram_cell[     428] = 32'h000000a9;
    ram_cell[     429] = 32'h0000011c;
    ram_cell[     430] = 32'h000001f3;
    ram_cell[     431] = 32'h0000006d;
    ram_cell[     432] = 32'h00000004;
    ram_cell[     433] = 32'h00000057;
    ram_cell[     434] = 32'h0000017e;
    ram_cell[     435] = 32'h00000126;
    ram_cell[     436] = 32'h0000013c;
    ram_cell[     437] = 32'h0000011d;
    ram_cell[     438] = 32'h00000086;
    ram_cell[     439] = 32'h000001ed;
    ram_cell[     440] = 32'h000000d5;
    ram_cell[     441] = 32'h000000ea;
    ram_cell[     442] = 32'h0000004b;
    ram_cell[     443] = 32'h00000136;
    ram_cell[     444] = 32'h000001a6;
    ram_cell[     445] = 32'h00000001;
    ram_cell[     446] = 32'h000001c9;
    ram_cell[     447] = 32'h000001e5;
    ram_cell[     448] = 32'h0000000b;
    ram_cell[     449] = 32'h000000b4;
    ram_cell[     450] = 32'h000001cc;
    ram_cell[     451] = 32'h000000bd;
    ram_cell[     452] = 32'h000001be;
    ram_cell[     453] = 32'h000001aa;
    ram_cell[     454] = 32'h0000012c;
    ram_cell[     455] = 32'h0000002c;
    ram_cell[     456] = 32'h000000c1;
    ram_cell[     457] = 32'h00000099;
    ram_cell[     458] = 32'h000001ba;
    ram_cell[     459] = 32'h00000041;
    ram_cell[     460] = 32'h00000183;
    ram_cell[     461] = 32'h000001bb;
    ram_cell[     462] = 32'h00000127;
    ram_cell[     463] = 32'h000001c4;
    ram_cell[     464] = 32'h000001d2;
    ram_cell[     465] = 32'h0000018b;
    ram_cell[     466] = 32'h00000177;
    ram_cell[     467] = 32'h00000079;
    ram_cell[     468] = 32'h0000016c;
    ram_cell[     469] = 32'h0000014e;
    ram_cell[     470] = 32'h00000040;
    ram_cell[     471] = 32'h000001ce;
    ram_cell[     472] = 32'h000001d5;
    ram_cell[     473] = 32'h000000a5;
    ram_cell[     474] = 32'h000000ee;
    ram_cell[     475] = 32'h000001fc;
    ram_cell[     476] = 32'h000000bf;
    ram_cell[     477] = 32'h00000142;
    ram_cell[     478] = 32'h000001f5;
    ram_cell[     479] = 32'h0000001e;
    ram_cell[     480] = 32'h00000090;
    ram_cell[     481] = 32'h00000184;
    ram_cell[     482] = 32'h0000014d;
    ram_cell[     483] = 32'h00000100;
    ram_cell[     484] = 32'h000000ad;
    ram_cell[     485] = 32'h00000051;
    ram_cell[     486] = 32'h00000002;
    ram_cell[     487] = 32'h00000174;
    ram_cell[     488] = 32'h000000e2;
    ram_cell[     489] = 32'h00000082;
    ram_cell[     490] = 32'h00000159;
    ram_cell[     491] = 32'h0000013b;
    ram_cell[     492] = 32'h0000002f;
    ram_cell[     493] = 32'h00000162;
    ram_cell[     494] = 32'h00000185;
    ram_cell[     495] = 32'h00000025;
    ram_cell[     496] = 32'h0000004a;
    ram_cell[     497] = 32'h000000c2;
    ram_cell[     498] = 32'h00000069;
    ram_cell[     499] = 32'h0000002e;
    ram_cell[     500] = 32'h000000e5;
    ram_cell[     501] = 32'h000000a1;
    ram_cell[     502] = 32'h00000124;
    ram_cell[     503] = 32'h00000046;
    ram_cell[     504] = 32'h00000150;
    ram_cell[     505] = 32'h00000135;
    ram_cell[     506] = 32'h00000137;
    ram_cell[     507] = 32'h0000017a;
    ram_cell[     508] = 32'h000001af;
    ram_cell[     509] = 32'h00000065;
    ram_cell[     510] = 32'h00000157;
    ram_cell[     511] = 32'h00000119;
end

endmodule

